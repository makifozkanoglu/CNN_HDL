`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/31/2020 03:30:08 PM
// Design Name: 
// Module Name: kernel_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module kernel_tb #(parameter BIT_SIZE = 9,
                   parameter INPUT_WIDTH=32,
                   parameter INPUT_HEIGHT=32,
                   parameter CHANNEL_SIZE=3, 
                   parameter SUBKERNEL_OUT_BIT = 24, //BIT_SIZE*2+ceil of log2(KERNEL_WIDTH*KERNEL_HEIGHT)
                   parameter KERNEL_WIDTH = 6, 
                   parameter KERNEL_HEIGHT = 6, 
                   parameter STRIDE = 1,
                   parameter OUTPUT_WIDTH = (INPUT_WIDTH - KERNEL_WIDTH) / STRIDE + 1,
                   parameter OUTPUT_HEIGHT = (INPUT_HEIGHT - KERNEL_HEIGHT) / STRIDE + 1,
                   parameter CHANNEL_EXTENSION_BIT = 2 //ceil of log2(CHANNEL_SIZE)
                   );
    
    wire [INPUT_WIDTH*INPUT_HEIGHT*CHANNEL_SIZE*BIT_SIZE-1:0] input_buffer;
    wire [KERNEL_WIDTH*KERNEL_HEIGHT*CHANNEL_SIZE*BIT_SIZE-1:0] kernel_buffer;
    wire [BIT_SIZE - 1:0] bias; assign bias=0;
    reg clock,reset,enable;
    wire [(SUBKERNEL_OUT_BIT + CHANNEL_EXTENSION_BIT)*OUTPUT_WIDTH*OUTPUT_HEIGHT - 1 :0] conv_result;
    
    genvar i,j,k;
    wire [SUBKERNEL_OUT_BIT + CHANNEL_EXTENSION_BIT - 1:0] conv_result_array_for_tb [OUTPUT_WIDTH-1:0][OUTPUT_HEIGHT-1:0]; //SUBKERNEL_OUT_BIT + 1 ==> ceil of log2(CHANNEL_SIZE)
    for (i=0;i<OUTPUT_HEIGHT;i=i+1) begin
        for (j=0;j<OUTPUT_WIDTH;j=j+1) begin
            assign conv_result_array_for_tb[j][i]=conv_result[(SUBKERNEL_OUT_BIT + 1)*(i*OUTPUT_WIDTH+j+1) - 1:(SUBKERNEL_OUT_BIT + 1)*(i*OUTPUT_WIDTH+j)];
        end
    end
    
    wire done;
    kernel #(BIT_SIZE,
             INPUT_WIDTH,
             INPUT_HEIGHT,
             CHANNEL_SIZE, 
             SUBKERNEL_OUT_BIT, 
             KERNEL_WIDTH, 
             KERNEL_HEIGHT, 
             STRIDE,
             OUTPUT_WIDTH,
             OUTPUT_HEIGHT,
             CHANNEL_EXTENSION_BIT)
           uut(input_buffer, 
               kernel_buffer,
               bias,
               clock,
               reset,
               enable,
               conv_result,
               done);
   
   
    reg [BIT_SIZE-1:0] input_array [INPUT_WIDTH-1:0][INPUT_HEIGHT-1:0][CHANNEL_SIZE-1:0];
    for (i=0;i<CHANNEL_SIZE;i=i+1) begin
        for (j=0;j<INPUT_HEIGHT;j=j+1) begin
            for (k=0;k<INPUT_WIDTH;k=k+1) begin
                assign input_buffer  [i*INPUT_WIDTH*INPUT_HEIGHT*BIT_SIZE+
                                     j*INPUT_WIDTH*BIT_SIZE+
                                     (k+1)*BIT_SIZE - 1:
                                     i*INPUT_WIDTH*INPUT_HEIGHT*BIT_SIZE+
                                     j*INPUT_WIDTH*BIT_SIZE+
                                     k*BIT_SIZE]=input_array[k][j][i];
            end
        end
    end
    
    
    reg [BIT_SIZE-1:0] kernel_array [KERNEL_WIDTH-1:0][KERNEL_HEIGHT-1:0][CHANNEL_SIZE-1:0];
    for (i=0;i<CHANNEL_SIZE;i=i+1) begin
        for (j=0;j<KERNEL_HEIGHT;j=j+1) begin
            for (k=0;k<KERNEL_WIDTH;k=k+1) begin
                assign kernel_buffer  [i*KERNEL_WIDTH*KERNEL_HEIGHT*BIT_SIZE+
                                      j*KERNEL_WIDTH*BIT_SIZE+
                                      (k+1)*BIT_SIZE - 1:
                                      i*KERNEL_WIDTH*KERNEL_HEIGHT*BIT_SIZE+
                                      j*KERNEL_WIDTH*BIT_SIZE+
                                      k*BIT_SIZE]=kernel_array[k][j][i];
            end
        end
    end
    integer a,b,c;
    reg [7:0] x;
    reg s;
    initial
    begin
        s=1;
        x=1;
        reset=1;
        clock=0;
        enable=0;
        #50;
        for (a=0;a<CHANNEL_SIZE;a=a+1) begin
            for (b=0;b<KERNEL_HEIGHT;b=b+1) begin
                for (c=0;c<KERNEL_WIDTH;c=c+1) begin
                    if(s)
                        kernel_array[c][b][a]=1;//8'd1;//x;//8'd1;
                    else
                        kernel_array[c][b][a]=-1;
                    s=~s;
                    //x=x+1;
                end
            end
        end
        for (a=0;a<CHANNEL_SIZE;a=a+1) begin
            for (b=0;b<INPUT_HEIGHT;b=b+1) begin
                for (c=0;c<INPUT_WIDTH;c=c+1) begin
                    input_array[c][b][a]=x;//8'd1;
                    x=x+1;
                end
            end
        end
        
        #20;
        reset=0;
        enable=1;
        
        wait (done);
        #20;
        reset=1;
        enable=0;
        #50;
        kernel_array[0][0][0]=95;
		kernel_array[1][0][0]=-16;
		kernel_array[2][0][0]=-89;
		kernel_array[3][0][0]=-29;
		kernel_array[4][0][0]=85;
		kernel_array[5][0][0]=-10;
		kernel_array[0][1][0]=-21;
		kernel_array[1][1][0]=52;
		kernel_array[2][1][0]=-70;
		kernel_array[3][1][0]=47;
		kernel_array[4][1][0]=100;
		kernel_array[5][1][0]=-21;
		kernel_array[0][2][0]=-31;
		kernel_array[1][2][0]=-7;
		kernel_array[2][2][0]=-89;
		kernel_array[3][2][0]=-28;
		kernel_array[4][2][0]=-58;
		kernel_array[5][2][0]=-29;
		kernel_array[0][3][0]=97;
		kernel_array[1][3][0]=5;
		kernel_array[2][3][0]=-61;
		kernel_array[3][3][0]=9;
		kernel_array[4][3][0]=69;
		kernel_array[5][3][0]=-43;
		kernel_array[0][4][0]=25;
		kernel_array[1][4][0]=65;
		kernel_array[2][4][0]=-89;
		kernel_array[3][4][0]=16;
		kernel_array[4][4][0]=-93;
		kernel_array[5][4][0]=-47;
		kernel_array[0][5][0]=48;
		kernel_array[1][5][0]=62;
		kernel_array[2][5][0]=0;
		kernel_array[3][5][0]=-36;
		kernel_array[4][5][0]=97;
		kernel_array[5][5][0]=77;
		kernel_array[0][0][1]=-47;
		kernel_array[1][0][1]=-96;
		kernel_array[2][0][1]=41;
		kernel_array[3][0][1]=-29;
		kernel_array[4][0][1]=24;
		kernel_array[5][0][1]=-66;
		kernel_array[0][1][1]=20;
		kernel_array[1][1][1]=-55;
		kernel_array[2][1][1]=-33;
		kernel_array[3][1][1]=-9;
		kernel_array[4][1][1]=-22;
		kernel_array[5][1][1]=-93;
		kernel_array[0][2][1]=-14;
		kernel_array[1][2][1]=18;
		kernel_array[2][2][1]=67;
		kernel_array[3][2][1]=-85;
		kernel_array[4][2][1]=-77;
		kernel_array[5][2][1]=62;
		kernel_array[0][3][1]=44;
		kernel_array[1][3][1]=86;
		kernel_array[2][3][1]=-15;
		kernel_array[3][3][1]=85;
		kernel_array[4][3][1]=103;
		kernel_array[5][3][1]=56;
		kernel_array[0][4][1]=-86;
		kernel_array[1][4][1]=78;
		kernel_array[2][4][1]=62;
		kernel_array[3][4][1]=-53;
		kernel_array[4][4][1]=-86;
		kernel_array[5][4][1]=-44;
		kernel_array[0][5][1]=0;
		kernel_array[1][5][1]=57;
		kernel_array[2][5][1]=42;
		kernel_array[3][5][1]=82;
		kernel_array[4][5][1]=-17;
		kernel_array[5][5][1]=24;
		kernel_array[0][0][2]=39;
		kernel_array[1][0][2]=13;
		kernel_array[2][0][2]=43;
		kernel_array[3][0][2]=18;
		kernel_array[4][0][2]=-23;
		kernel_array[5][0][2]=-65;
		kernel_array[0][1][2]=-64;
		kernel_array[1][1][2]=-63;
		kernel_array[2][1][2]=78;
		kernel_array[3][1][2]=-64;
		kernel_array[4][1][2]=-87;
		kernel_array[5][1][2]=76;
		kernel_array[0][2][2]=-92;
		kernel_array[1][2][2]=-16;
		kernel_array[2][2][2]=0;
		kernel_array[3][2][2]=9;
		kernel_array[4][2][2]=-31;
		kernel_array[5][2][2]=-48;
		kernel_array[0][3][2]=-91;
		kernel_array[1][3][2]=97;
		kernel_array[2][3][2]=-94;
		kernel_array[3][3][2]=26;
		kernel_array[4][3][2]=-17;
		kernel_array[5][3][2]=26;
		kernel_array[0][4][2]=89;
		kernel_array[1][4][2]=32;
		kernel_array[2][4][2]=-88;
		kernel_array[3][4][2]=-33;
		kernel_array[4][4][2]=96;
		kernel_array[5][4][2]=10;
		kernel_array[0][5][2]=34;
		kernel_array[1][5][2]=-34;
		kernel_array[2][5][2]=-72;
		kernel_array[3][5][2]=-9;
		kernel_array[4][5][2]=-48;
		kernel_array[5][5][2]=-58;
        
        /*
        
        
        sdadas
        */
        
        input_array[0][0][0]=28;
		input_array[1][0][0]=37;
		input_array[2][0][0]=38;
		input_array[3][0][0]=42;
		input_array[4][0][0]=44;
		input_array[5][0][0]=40;
		input_array[6][0][0]=40;
		input_array[7][0][0]=24;
		input_array[8][0][0]=32;
		input_array[9][0][0]=43;
		input_array[10][0][0]=30;
		input_array[11][0][0]=32;
		input_array[12][0][0]=41;
		input_array[13][0][0]=52;
		input_array[14][0][0]=67;
		input_array[15][0][0]=50;
		input_array[16][0][0]=44;
		input_array[17][0][0]=43;
		input_array[18][0][0]=38;
		input_array[19][0][0]=38;
		input_array[20][0][0]=41;
		input_array[21][0][0]=47;
		input_array[22][0][0]=62;
		input_array[23][0][0]=87;
		input_array[24][0][0]=60;
		input_array[25][0][0]=49;
		input_array[26][0][0]=63;
		input_array[27][0][0]=59;
		input_array[28][0][0]=48;
		input_array[29][0][0]=76;
		input_array[30][0][0]=81;
		input_array[31][0][0]=85;
		input_array[0][1][0]=33;
		input_array[1][1][0]=34;
		input_array[2][1][0]=32;
		input_array[3][1][0]=39;
		input_array[4][1][0]=35;
		input_array[5][1][0]=38;
		input_array[6][1][0]=38;
		input_array[7][1][0]=40;
		input_array[8][1][0]=54;
		input_array[9][1][0]=48;
		input_array[10][1][0]=28;
		input_array[11][1][0]=40;
		input_array[12][1][0]=56;
		input_array[13][1][0]=66;
		input_array[14][1][0]=79;
		input_array[15][1][0]=47;
		input_array[16][1][0]=42;
		input_array[17][1][0]=50;
		input_array[18][1][0]=64;
		input_array[19][1][0]=47;
		input_array[20][1][0]=55;
		input_array[21][1][0]=81;
		input_array[22][1][0]=84;
		input_array[23][1][0]=109;
		input_array[24][1][0]=92;
		input_array[25][1][0]=59;
		input_array[26][1][0]=69;
		input_array[27][1][0]=79;
		input_array[28][1][0]=71;
		input_array[29][1][0]=95;
		input_array[30][1][0]=96;
		input_array[31][1][0]=85;
		input_array[0][2][0]=39;
		input_array[1][2][0]=40;
		input_array[2][2][0]=57;
		input_array[3][2][0]=46;
		input_array[4][2][0]=44;
		input_array[5][2][0]=40;
		input_array[6][2][0]=41;
		input_array[7][2][0]=66;
		input_array[8][2][0]=90;
		input_array[9][2][0]=57;
		input_array[10][2][0]=48;
		input_array[11][2][0]=72;
		input_array[12][2][0]=74;
		input_array[13][2][0]=76;
		input_array[14][2][0]=93;
		input_array[15][2][0]=66;
		input_array[16][2][0]=65;
		input_array[17][2][0]=80;
		input_array[18][2][0]=90;
		input_array[19][2][0]=67;
		input_array[20][2][0]=88;
		input_array[21][2][0]=96;
		input_array[22][2][0]=83;
		input_array[23][2][0]=105;
		input_array[24][2][0]=107;
		input_array[25][2][0]=86;
		input_array[26][2][0]=89;
		input_array[27][2][0]=93;
		input_array[28][2][0]=86;
		input_array[29][2][0]=93;
		input_array[30][2][0]=107;
		input_array[31][2][0]=95;
		input_array[0][3][0]=54;
		input_array[1][3][0]=62;
		input_array[2][3][0]=84;
		input_array[3][3][0]=62;
		input_array[4][3][0]=70;
		input_array[5][3][0]=55;
		input_array[6][3][0]=78;
		input_array[7][3][0]=85;
		input_array[8][3][0]=99;
		input_array[9][3][0]=84;
		input_array[10][3][0]=95;
		input_array[11][3][0]=90;
		input_array[12][3][0]=96;
		input_array[13][3][0]=103;
		input_array[14][3][0]=93;
		input_array[15][3][0]=95;
		input_array[16][3][0]=94;
		input_array[17][3][0]=100;
		input_array[18][3][0]=94;
		input_array[19][3][0]=87;
		input_array[20][3][0]=92;
		input_array[21][3][0]=89;
		input_array[22][3][0]=96;
		input_array[23][3][0]=96;
		input_array[24][3][0]=83;
		input_array[25][3][0]=76;
		input_array[26][3][0]=95;
		input_array[27][3][0]=104;
		input_array[28][3][0]=97;
		input_array[29][3][0]=101;
		input_array[30][3][0]=99;
		input_array[31][3][0]=91;
		input_array[0][4][0]=74;
		input_array[1][4][0]=72;
		input_array[2][4][0]=78;
		input_array[3][4][0]=85;
		input_array[4][4][0]=95;
		input_array[5][4][0]=77;
		input_array[6][4][0]=103;
		input_array[7][4][0]=98;
		input_array[8][4][0]=80;
		input_array[9][4][0]=93;
		input_array[10][4][0]=99;
		input_array[11][4][0]=93;
		input_array[12][4][0]=101;
		input_array[13][4][0]=105;
		input_array[14][4][0]=84;
		input_array[15][4][0]=84;
		input_array[16][4][0]=86;
		input_array[17][4][0]=87;
		input_array[18][4][0]=80;
		input_array[19][4][0]=87;
		input_array[20][4][0]=80;
		input_array[21][4][0]=91;
		input_array[22][4][0]=93;
		input_array[23][4][0]=74;
		input_array[24][4][0]=81;
		input_array[25][4][0]=77;
		input_array[26][4][0]=89;
		input_array[27][4][0]=82;
		input_array[28][4][0]=84;
		input_array[29][4][0]=78;
		input_array[30][4][0]=72;
		input_array[31][4][0]=84;
		input_array[0][5][0]=76;
		input_array[1][5][0]=68;
		input_array[2][5][0]=69;
		input_array[3][5][0]=74;
		input_array[4][5][0]=78;
		input_array[5][5][0]=81;
		input_array[6][5][0]=89;
		input_array[7][5][0]=90;
		input_array[8][5][0]=79;
		input_array[9][5][0]=66;
		input_array[10][5][0]=81;
		input_array[11][5][0]=91;
		input_array[12][5][0]=87;
		input_array[13][5][0]=86;
		input_array[14][5][0]=90;
		input_array[15][5][0]=85;
		input_array[16][5][0]=81;
		input_array[17][5][0]=82;
		input_array[18][5][0]=78;
		input_array[19][5][0]=85;
		input_array[20][5][0]=87;
		input_array[21][5][0]=91;
		input_array[22][5][0]=83;
		input_array[23][5][0]=80;
		input_array[24][5][0]=87;
		input_array[25][5][0]=91;
		input_array[26][5][0]=98;
		input_array[27][5][0]=74;
		input_array[28][5][0]=59;
		input_array[29][5][0]=71;
		input_array[30][5][0]=72;
		input_array[31][5][0]=94;
		input_array[0][6][0]=77;
		input_array[1][6][0]=74;
		input_array[2][6][0]=73;
		input_array[3][6][0]=70;
		input_array[4][6][0]=67;
		input_array[5][6][0]=84;
		input_array[6][6][0]=94;
		input_array[7][6][0]=98;
		input_array[8][6][0]=82;
		input_array[9][6][0]=72;
		input_array[10][6][0]=75;
		input_array[11][6][0]=75;
		input_array[12][6][0]=81;
		input_array[13][6][0]=87;
		input_array[14][6][0]=91;
		input_array[15][6][0]=82;
		input_array[16][6][0]=90;
		input_array[17][6][0]=85;
		input_array[18][6][0]=95;
		input_array[19][6][0]=103;
		input_array[20][6][0]=104;
		input_array[21][6][0]=91;
		input_array[22][6][0]=78;
		input_array[23][6][0]=79;
		input_array[24][6][0]=95;
		input_array[25][6][0]=95;
		input_array[26][6][0]=91;
		input_array[27][6][0]=71;
		input_array[28][6][0]=65;
		input_array[29][6][0]=85;
		input_array[30][6][0]=80;
		input_array[31][6][0]=80;
		input_array[0][7][0]=79;
		input_array[1][7][0]=76;
		input_array[2][7][0]=85;
		input_array[3][7][0]=77;
		input_array[4][7][0]=83;
		input_array[5][7][0]=81;
		input_array[6][7][0]=94;
		input_array[7][7][0]=122;
		input_array[8][7][0]=94;
		input_array[9][7][0]=82;
		input_array[10][7][0]=93;
		input_array[11][7][0]=86;
		input_array[12][7][0]=101;
		input_array[13][7][0]=91;
		input_array[14][7][0]=91;
		input_array[15][7][0]=102;
		input_array[16][7][0]=95;
		input_array[17][7][0]=93;
		input_array[18][7][0]=100;
		input_array[19][7][0]=111;
		input_array[20][7][0]=103;
		input_array[21][7][0]=98;
		input_array[22][7][0]=93;
		input_array[23][7][0]=78;
		input_array[24][7][0]=90;
		input_array[25][7][0]=93;
		input_array[26][7][0]=83;
		input_array[27][7][0]=71;
		input_array[28][7][0]=74;
		input_array[29][7][0]=89;
		input_array[30][7][0]=77;
		input_array[31][7][0]=56;
		input_array[0][8][0]=52;
		input_array[1][8][0]=51;
		input_array[2][8][0]=62;
		input_array[3][8][0]=74;
		input_array[4][8][0]=75;
		input_array[5][8][0]=87;
		input_array[6][8][0]=121;
		input_array[7][8][0]=129;
		input_array[8][8][0]=97;
		input_array[9][8][0]=99;
		input_array[10][8][0]=115;
		input_array[11][8][0]=128;
		input_array[12][8][0]=121;
		input_array[13][8][0]=83;
		input_array[14][8][0]=99;
		input_array[15][8][0]=95;
		input_array[16][8][0]=87;
		input_array[17][8][0]=92;
		input_array[18][8][0]=95;
		input_array[19][8][0]=103;
		input_array[20][8][0]=101;
		input_array[21][8][0]=101;
		input_array[22][8][0]=86;
		input_array[23][8][0]=74;
		input_array[24][8][0]=84;
		input_array[25][8][0]=105;
		input_array[26][8][0]=111;
		input_array[27][8][0]=74;
		input_array[28][8][0]=93;
		input_array[29][8][0]=94;
		input_array[30][8][0]=91;
		input_array[31][8][0]=75;
		input_array[0][9][0]=45;
		input_array[1][9][0]=27;
		input_array[2][9][0]=37;
		input_array[3][9][0]=55;
		input_array[4][9][0]=60;
		input_array[5][9][0]=83;
		input_array[6][9][0]=113;
		input_array[7][9][0]=109;
		input_array[8][9][0]=97;
		input_array[9][9][0]=102;
		input_array[10][9][0]=108;
		input_array[11][9][0]=136;
		input_array[12][9][0]=89;
		input_array[13][9][0]=95;
		input_array[14][9][0]=111;
		input_array[15][9][0]=104;
		input_array[16][9][0]=112;
		input_array[17][9][0]=113;
		input_array[18][9][0]=109;
		input_array[19][9][0]=117;
		input_array[20][9][0]=104;
		input_array[21][9][0]=111;
		input_array[22][9][0]=77;
		input_array[23][9][0]=74;
		input_array[24][9][0]=96;
		input_array[25][9][0]=97;
		input_array[26][9][0]=101;
		input_array[27][9][0]=83;
		input_array[28][9][0]=106;
		input_array[29][9][0]=88;
		input_array[30][9][0]=80;
		input_array[31][9][0]=88;
		input_array[0][10][0]=67;
		input_array[1][10][0]=41;
		input_array[2][10][0]=54;
		input_array[3][10][0]=54;
		input_array[4][10][0]=63;
		input_array[5][10][0]=92;
		input_array[6][10][0]=112;
		input_array[7][10][0]=99;
		input_array[8][10][0]=91;
		input_array[9][10][0]=104;
		input_array[10][10][0]=149;
		input_array[11][10][0]=125;
		input_array[12][10][0]=82;
		input_array[13][10][0]=109;
		input_array[14][10][0]=107;
		input_array[15][10][0]=102;
		input_array[16][10][0]=122;
		input_array[17][10][0]=116;
		input_array[18][10][0]=116;
		input_array[19][10][0]=120;
		input_array[20][10][0]=93;
		input_array[21][10][0]=89;
		input_array[22][10][0]=92;
		input_array[23][10][0]=80;
		input_array[24][10][0]=93;
		input_array[25][10][0]=100;
		input_array[26][10][0]=96;
		input_array[27][10][0]=110;
		input_array[28][10][0]=108;
		input_array[29][10][0]=71;
		input_array[30][10][0]=69;
		input_array[31][10][0]=96;
		input_array[0][11][0]=79;
		input_array[1][11][0]=82;
		input_array[2][11][0]=91;
		input_array[3][11][0]=93;
		input_array[4][11][0]=69;
		input_array[5][11][0]=88;
		input_array[6][11][0]=123;
		input_array[7][11][0]=96;
		input_array[8][11][0]=94;
		input_array[9][11][0]=105;
		input_array[10][11][0]=136;
		input_array[11][11][0]=104;
		input_array[12][11][0]=77;
		input_array[13][11][0]=109;
		input_array[14][11][0]=95;
		input_array[15][11][0]=93;
		input_array[16][11][0]=112;
		input_array[17][11][0]=100;
		input_array[18][11][0]=114;
		input_array[19][11][0]=114;
		input_array[20][11][0]=92;
		input_array[21][11][0]=92;
		input_array[22][11][0]=106;
		input_array[23][11][0]=101;
		input_array[24][11][0]=105;
		input_array[25][11][0]=118;
		input_array[26][11][0]=121;
		input_array[27][11][0]=119;
		input_array[28][11][0]=86;
		input_array[29][11][0]=72;
		input_array[30][11][0]=75;
		input_array[31][11][0]=83;
		input_array[0][12][0]=91;
		input_array[1][12][0]=102;
		input_array[2][12][0]=107;
		input_array[3][12][0]=122;
		input_array[4][12][0]=102;
		input_array[5][12][0]=85;
		input_array[6][12][0]=80;
		input_array[7][12][0]=76;
		input_array[8][12][0]=83;
		input_array[9][12][0]=112;
		input_array[10][12][0]=110;
		input_array[11][12][0]=85;
		input_array[12][12][0]=69;
		input_array[13][12][0]=95;
		input_array[14][12][0]=95;
		input_array[15][12][0]=92;
		input_array[16][12][0]=96;
		input_array[17][12][0]=91;
		input_array[18][12][0]=94;
		input_array[19][12][0]=104;
		input_array[20][12][0]=110;
		input_array[21][12][0]=111;
		input_array[22][12][0]=104;
		input_array[23][12][0]=100;
		input_array[24][12][0]=96;
		input_array[25][12][0]=104;
		input_array[26][12][0]=100;
		input_array[27][12][0]=93;
		input_array[28][12][0]=83;
		input_array[29][12][0]=81;
		input_array[30][12][0]=81;
		input_array[31][12][0]=87;
		input_array[0][13][0]=119;
		input_array[1][13][0]=116;
		input_array[2][13][0]=133;
		input_array[3][13][0]=136;
		input_array[4][13][0]=127;
		input_array[5][13][0]=126;
		input_array[6][13][0]=59;
		input_array[7][13][0]=57;
		input_array[8][13][0]=73;
		input_array[9][13][0]=88;
		input_array[10][13][0]=111;
		input_array[11][13][0]=101;
		input_array[12][13][0]=69;
		input_array[13][13][0]=75;
		input_array[14][13][0]=91;
		input_array[15][13][0]=102;
		input_array[16][13][0]=117;
		input_array[17][13][0]=130;
		input_array[18][13][0]=143;
		input_array[19][13][0]=154;
		input_array[20][13][0]=150;
		input_array[21][13][0]=116;
		input_array[22][13][0]=114;
		input_array[23][13][0]=104;
		input_array[24][13][0]=94;
		input_array[25][13][0]=98;
		input_array[26][13][0]=101;
		input_array[27][13][0]=94;
		input_array[28][13][0]=92;
		input_array[29][13][0]=89;
		input_array[30][13][0]=84;
		input_array[31][13][0]=82;
		input_array[0][14][0]=118;
		input_array[1][14][0]=123;
		input_array[2][14][0]=136;
		input_array[3][14][0]=131;
		input_array[4][14][0]=134;
		input_array[5][14][0]=133;
		input_array[6][14][0]=56;
		input_array[7][14][0]=58;
		input_array[8][14][0]=75;
		input_array[9][14][0]=88;
		input_array[10][14][0]=142;
		input_array[11][14][0]=162;
		input_array[12][14][0]=129;
		input_array[13][14][0]=136;
		input_array[14][14][0]=150;
		input_array[15][14][0]=153;
		input_array[16][14][0]=131;
		input_array[17][14][0]=189;
		input_array[18][14][0]=213;
		input_array[19][14][0]=209;
		input_array[20][14][0]=195;
		input_array[21][14][0]=133;
		input_array[22][14][0]=114;
		input_array[23][14][0]=108;
		input_array[24][14][0]=115;
		input_array[25][14][0]=113;
		input_array[26][14][0]=111;
		input_array[27][14][0]=116;
		input_array[28][14][0]=99;
		input_array[29][14][0]=98;
		input_array[30][14][0]=83;
		input_array[31][14][0]=79;
		input_array[0][15][0]=88;
		input_array[1][15][0]=100;
		input_array[2][15][0]=110;
		input_array[3][15][0]=126;
		input_array[4][15][0]=125;
		input_array[5][15][0]=122;
		input_array[6][15][0]=66;
		input_array[7][15][0]=60;
		input_array[8][15][0]=97;
		input_array[9][15][0]=104;
		input_array[10][15][0]=177;
		input_array[11][15][0]=184;
		input_array[12][15][0]=164;
		input_array[13][15][0]=170;
		input_array[14][15][0]=179;
		input_array[15][15][0]=181;
		input_array[16][15][0]=152;
		input_array[17][15][0]=182;
		input_array[18][15][0]=208;
		input_array[19][15][0]=227;
		input_array[20][15][0]=211;
		input_array[21][15][0]=164;
		input_array[22][15][0]=140;
		input_array[23][15][0]=126;
		input_array[24][15][0]=132;
		input_array[25][15][0]=136;
		input_array[26][15][0]=132;
		input_array[27][15][0]=135;
		input_array[28][15][0]=113;
		input_array[29][15][0]=116;
		input_array[30][15][0]=97;
		input_array[31][15][0]=109;
		input_array[0][16][0]=78;
		input_array[1][16][0]=86;
		input_array[2][16][0]=94;
		input_array[3][16][0]=128;
		input_array[4][16][0]=126;
		input_array[5][16][0]=114;
		input_array[6][16][0]=95;
		input_array[7][16][0]=53;
		input_array[8][16][0]=102;
		input_array[9][16][0]=129;
		input_array[10][16][0]=198;
		input_array[11][16][0]=201;
		input_array[12][16][0]=189;
		input_array[13][16][0]=195;
		input_array[14][16][0]=205;
		input_array[15][16][0]=208;
		input_array[16][16][0]=181;
		input_array[17][16][0]=173;
		input_array[18][16][0]=190;
		input_array[19][16][0]=207;
		input_array[20][16][0]=216;
		input_array[21][16][0]=174;
		input_array[22][16][0]=154;
		input_array[23][16][0]=126;
		input_array[24][16][0]=131;
		input_array[25][16][0]=145;
		input_array[26][16][0]=146;
		input_array[27][16][0]=141;
		input_array[28][16][0]=127;
		input_array[29][16][0]=124;
		input_array[30][16][0]=111;
		input_array[31][16][0]=116;
		input_array[0][17][0]=80;
		input_array[1][17][0]=79;
		input_array[2][17][0]=93;
		input_array[3][17][0]=121;
		input_array[4][17][0]=128;
		input_array[5][17][0]=116;
		input_array[6][17][0]=92;
		input_array[7][17][0]=40;
		input_array[8][17][0]=92;
		input_array[9][17][0]=162;
		input_array[10][17][0]=207;
		input_array[11][17][0]=219;
		input_array[12][17][0]=216;
		input_array[13][17][0]=211;
		input_array[14][17][0]=208;
		input_array[15][17][0]=211;
		input_array[16][17][0]=201;
		input_array[17][17][0]=179;
		input_array[18][17][0]=165;
		input_array[19][17][0]=139;
		input_array[20][17][0]=175;
		input_array[21][17][0]=152;
		input_array[22][17][0]=126;
		input_array[23][17][0]=122;
		input_array[24][17][0]=142;
		input_array[25][17][0]=150;
		input_array[26][17][0]=157;
		input_array[27][17][0]=153;
		input_array[28][17][0]=134;
		input_array[29][17][0]=132;
		input_array[30][17][0]=134;
		input_array[31][17][0]=120;
		input_array[0][18][0]=104;
		input_array[1][18][0]=111;
		input_array[2][18][0]=121;
		input_array[3][18][0]=130;
		input_array[4][18][0]=126;
		input_array[5][18][0]=121;
		input_array[6][18][0]=106;
		input_array[7][18][0]=75;
		input_array[8][18][0]=108;
		input_array[9][18][0]=188;
		input_array[10][18][0]=219;
		input_array[11][18][0]=233;
		input_array[12][18][0]=225;
		input_array[13][18][0]=222;
		input_array[14][18][0]=208;
		input_array[15][18][0]=219;
		input_array[16][18][0]=216;
		input_array[17][18][0]=177;
		input_array[18][18][0]=136;
		input_array[19][18][0]=97;
		input_array[20][18][0]=115;
		input_array[21][18][0]=101;
		input_array[22][18][0]=96;
		input_array[23][18][0]=138;
		input_array[24][18][0]=154;
		input_array[25][18][0]=151;
		input_array[26][18][0]=157;
		input_array[27][18][0]=152;
		input_array[28][18][0]=142;
		input_array[29][18][0]=139;
		input_array[30][18][0]=140;
		input_array[31][18][0]=116;
		input_array[0][19][0]=103;
		input_array[1][19][0]=119;
		input_array[2][19][0]=126;
		input_array[3][19][0]=135;
		input_array[4][19][0]=122;
		input_array[5][19][0]=116;
		input_array[6][19][0]=121;
		input_array[7][19][0]=123;
		input_array[8][19][0]=132;
		input_array[9][19][0]=193;
		input_array[10][19][0]=223;
		input_array[11][19][0]=230;
		input_array[12][19][0]=225;
		input_array[13][19][0]=229;
		input_array[14][19][0]=220;
		input_array[15][19][0]=226;
		input_array[16][19][0]=225;
		input_array[17][19][0]=182;
		input_array[18][19][0]=94;
		input_array[19][19][0]=83;
		input_array[20][19][0]=97;
		input_array[21][19][0]=90;
		input_array[22][19][0]=96;
		input_array[23][19][0]=140;
		input_array[24][19][0]=153;
		input_array[25][19][0]=149;
		input_array[26][19][0]=143;
		input_array[27][19][0]=130;
		input_array[28][19][0]=134;
		input_array[29][19][0]=128;
		input_array[30][19][0]=124;
		input_array[31][19][0]=110;
		input_array[0][20][0]=97;
		input_array[1][20][0]=106;
		input_array[2][20][0]=121;
		input_array[3][20][0]=117;
		input_array[4][20][0]=112;
		input_array[5][20][0]=122;
		input_array[6][20][0]=125;
		input_array[7][20][0]=109;
		input_array[8][20][0]=116;
		input_array[9][20][0]=178;
		input_array[10][20][0]=218;
		input_array[11][20][0]=222;
		input_array[12][20][0]=227;
		input_array[13][20][0]=234;
		input_array[14][20][0]=219;
		input_array[15][20][0]=226;
		input_array[16][20][0]=219;
		input_array[17][20][0]=192;
		input_array[18][20][0]=70;
		input_array[19][20][0]=63;
		input_array[20][20][0]=76;
		input_array[21][20][0]=82;
		input_array[22][20][0]=93;
		input_array[23][20][0]=130;
		input_array[24][20][0]=136;
		input_array[25][20][0]=143;
		input_array[26][20][0]=128;
		input_array[27][20][0]=104;
		input_array[28][20][0]=103;
		input_array[29][20][0]=103;
		input_array[30][20][0]=104;
		input_array[31][20][0]=113;
		input_array[0][21][0]=77;
		input_array[1][21][0]=103;
		input_array[2][21][0]=108;
		input_array[3][21][0]=104;
		input_array[4][21][0]=122;
		input_array[5][21][0]=109;
		input_array[6][21][0]=105;
		input_array[7][21][0]=98;
		input_array[8][21][0]=107;
		input_array[9][21][0]=138;
		input_array[10][21][0]=180;
		input_array[11][21][0]=186;
		input_array[12][21][0]=216;
		input_array[13][21][0]=229;
		input_array[14][21][0]=211;
		input_array[15][21][0]=216;
		input_array[16][21][0]=212;
		input_array[17][21][0]=199;
		input_array[18][21][0]=54;
		input_array[19][21][0]=16;
		input_array[20][21][0]=49;
		input_array[21][21][0]=67;
		input_array[22][21][0]=86;
		input_array[23][21][0]=119;
		input_array[24][21][0]=113;
		input_array[25][21][0]=117;
		input_array[26][21][0]=104;
		input_array[27][21][0]=87;
		input_array[28][21][0]=85;
		input_array[29][21][0]=86;
		input_array[30][21][0]=91;
		input_array[31][21][0]=93;
		input_array[0][22][0]=48;
		input_array[1][22][0]=82;
		input_array[2][22][0]=78;
		input_array[3][22][0]=107;
		input_array[4][22][0]=111;
		input_array[5][22][0]=95;
		input_array[6][22][0]=91;
		input_array[7][22][0]=94;
		input_array[8][22][0]=97;
		input_array[9][22][0]=97;
		input_array[10][22][0]=142;
		input_array[11][22][0]=116;
		input_array[12][22][0]=136;
		input_array[13][22][0]=151;
		input_array[14][22][0]=114;
		input_array[15][22][0]=113;
		input_array[16][22][0]=191;
		input_array[17][22][0]=198;
		input_array[18][22][0]=71;
		input_array[19][22][0]=25;
		input_array[20][22][0]=30;
		input_array[21][22][0]=47;
		input_array[22][22][0]=72;
		input_array[23][22][0]=105;
		input_array[24][22][0]=94;
		input_array[25][22][0]=84;
		input_array[26][22][0]=86;
		input_array[27][22][0]=78;
		input_array[28][22][0]=79;
		input_array[29][22][0]=77;
		input_array[30][22][0]=69;
		input_array[31][22][0]=89;
		input_array[0][23][0]=44;
		input_array[1][23][0]=63;
		input_array[2][23][0]=77;
		input_array[3][23][0]=93;
		input_array[4][23][0]=96;
		input_array[5][23][0]=93;
		input_array[6][23][0]=80;
		input_array[7][23][0]=82;
		input_array[8][23][0]=81;
		input_array[9][23][0]=94;
		input_array[10][23][0]=120;
		input_array[11][23][0]=68;
		input_array[12][23][0]=79;
		input_array[13][23][0]=72;
		input_array[14][23][0]=72;
		input_array[15][23][0]=78;
		input_array[16][23][0]=150;
		input_array[17][23][0]=173;
		input_array[18][23][0]=84;
		input_array[19][23][0]=49;
		input_array[20][23][0]=30;
		input_array[21][23][0]=48;
		input_array[22][23][0]=50;
		input_array[23][23][0]=100;
		input_array[24][23][0]=91;
		input_array[25][23][0]=77;
		input_array[26][23][0]=67;
		input_array[27][23][0]=63;
		input_array[28][23][0]=60;
		input_array[29][23][0]=73;
		input_array[30][23][0]=63;
		input_array[31][23][0]=78;
		input_array[0][24][0]=61;
		input_array[1][24][0]=77;
		input_array[2][24][0]=85;
		input_array[3][24][0]=75;
		input_array[4][24][0]=84;
		input_array[5][24][0]=79;
		input_array[6][24][0]=73;
		input_array[7][24][0]=77;
		input_array[8][24][0]=83;
		input_array[9][24][0]=88;
		input_array[10][24][0]=98;
		input_array[11][24][0]=60;
		input_array[12][24][0]=86;
		input_array[13][24][0]=107;
		input_array[14][24][0]=102;
		input_array[15][24][0]=88;
		input_array[16][24][0]=118;
		input_array[17][24][0]=156;
		input_array[18][24][0]=86;
		input_array[19][24][0]=61;
		input_array[20][24][0]=50;
		input_array[21][24][0]=64;
		input_array[22][24][0]=52;
		input_array[23][24][0]=68;
		input_array[24][24][0]=103;
		input_array[25][24][0]=85;
		input_array[26][24][0]=71;
		input_array[27][24][0]=67;
		input_array[28][24][0]=53;
		input_array[29][24][0]=90;
		input_array[30][24][0]=82;
		input_array[31][24][0]=75;
		input_array[0][25][0]=48;
		input_array[1][25][0]=59;
		input_array[2][25][0]=85;
		input_array[3][25][0]=81;
		input_array[4][25][0]=74;
		input_array[5][25][0]=85;
		input_array[6][25][0]=80;
		input_array[7][25][0]=81;
		input_array[8][25][0]=88;
		input_array[9][25][0]=89;
		input_array[10][25][0]=88;
		input_array[11][25][0]=66;
		input_array[12][25][0]=98;
		input_array[13][25][0]=102;
		input_array[14][25][0]=98;
		input_array[15][25][0]=96;
		input_array[16][25][0]=116;
		input_array[17][25][0]=143;
		input_array[18][25][0]=123;
		input_array[19][25][0]=82;
		input_array[20][25][0]=57;
		input_array[21][25][0]=49;
		input_array[22][25][0]=86;
		input_array[23][25][0]=58;
		input_array[24][25][0]=98;
		input_array[25][25][0]=86;
		input_array[26][25][0]=59;
		input_array[27][25][0]=57;
		input_array[28][25][0]=65;
		input_array[29][25][0]=102;
		input_array[30][25][0]=79;
		input_array[31][25][0]=78;
		input_array[0][26][0]=58;
		input_array[1][26][0]=56;
		input_array[2][26][0]=78;
		input_array[3][26][0]=82;
		input_array[4][26][0]=79;
		input_array[5][26][0]=88;
		input_array[6][26][0]=85;
		input_array[7][26][0]=87;
		input_array[8][26][0]=92;
		input_array[9][26][0]=92;
		input_array[10][26][0]=85;
		input_array[11][26][0]=67;
		input_array[12][26][0]=108;
		input_array[13][26][0]=95;
		input_array[14][26][0]=104;
		input_array[15][26][0]=83;
		input_array[16][26][0]=100;
		input_array[17][26][0]=133;
		input_array[18][26][0]=133;
		input_array[19][26][0]=94;
		input_array[20][26][0]=80;
		input_array[21][26][0]=60;
		input_array[22][26][0]=96;
		input_array[23][26][0]=80;
		input_array[24][26][0]=85;
		input_array[25][26][0]=79;
		input_array[26][26][0]=61;
		input_array[27][26][0]=73;
		input_array[28][26][0]=86;
		input_array[29][26][0]=88;
		input_array[30][26][0]=59;
		input_array[31][26][0]=58;
		input_array[0][27][0]=66;
		input_array[1][27][0]=68;
		input_array[2][27][0]=69;
		input_array[3][27][0]=76;
		input_array[4][27][0]=85;
		input_array[5][27][0]=89;
		input_array[6][27][0]=91;
		input_array[7][27][0]=91;
		input_array[8][27][0]=106;
		input_array[9][27][0]=98;
		input_array[10][27][0]=86;
		input_array[11][27][0]=71;
		input_array[12][27][0]=99;
		input_array[13][27][0]=98;
		input_array[14][27][0]=99;
		input_array[15][27][0]=77;
		input_array[16][27][0]=75;
		input_array[17][27][0]=118;
		input_array[18][27][0]=113;
		input_array[19][27][0]=103;
		input_array[20][27][0]=102;
		input_array[21][27][0]=101;
		input_array[22][27][0]=81;
		input_array[23][27][0]=98;
		input_array[24][27][0]=98;
		input_array[25][27][0]=86;
		input_array[26][27][0]=100;
		input_array[27][27][0]=98;
		input_array[28][27][0]=88;
		input_array[29][27][0]=78;
		input_array[30][27][0]=77;
		input_array[31][27][0]=72;
		input_array[0][28][0]=72;
		input_array[1][28][0]=82;
		input_array[2][28][0]=79;
		input_array[3][28][0]=82;
		input_array[4][28][0]=88;
		input_array[5][28][0]=86;
		input_array[6][28][0]=85;
		input_array[7][28][0]=84;
		input_array[8][28][0]=93;
		input_array[9][28][0]=84;
		input_array[10][28][0]=87;
		input_array[11][28][0]=79;
		input_array[12][28][0]=93;
		input_array[13][28][0]=88;
		input_array[14][28][0]=78;
		input_array[15][28][0]=83;
		input_array[16][28][0]=96;
		input_array[17][28][0]=118;
		input_array[18][28][0]=108;
		input_array[19][28][0]=106;
		input_array[20][28][0]=112;
		input_array[21][28][0]=111;
		input_array[22][28][0]=94;
		input_array[23][28][0]=105;
		input_array[24][28][0]=121;
		input_array[25][28][0]=97;
		input_array[26][28][0]=101;
		input_array[27][28][0]=90;
		input_array[28][28][0]=79;
		input_array[29][28][0]=86;
		input_array[30][28][0]=87;
		input_array[31][28][0]=87;
		input_array[0][29][0]=83;
		input_array[1][29][0]=87;
		input_array[2][29][0]=84;
		input_array[3][29][0]=92;
		input_array[4][29][0]=80;
		input_array[5][29][0]=83;
		input_array[6][29][0]=89;
		input_array[7][29][0]=98;
		input_array[8][29][0]=104;
		input_array[9][29][0]=102;
		input_array[10][29][0]=93;
		input_array[11][29][0]=110;
		input_array[12][29][0]=102;
		input_array[13][29][0]=109;
		input_array[14][29][0]=114;
		input_array[15][29][0]=113;
		input_array[16][29][0]=108;
		input_array[17][29][0]=114;
		input_array[18][29][0]=117;
		input_array[19][29][0]=122;
		input_array[20][29][0]=122;
		input_array[21][29][0]=117;
		input_array[22][29][0]=114;
		input_array[23][29][0]=120;
		input_array[24][29][0]=124;
		input_array[25][29][0]=104;
		input_array[26][29][0]=103;
		input_array[27][29][0]=100;
		input_array[28][29][0]=99;
		input_array[29][29][0]=99;
		input_array[30][29][0]=90;
		input_array[31][29][0]=81;
		input_array[0][30][0]=88;
		input_array[1][30][0]=90;
		input_array[2][30][0]=93;
		input_array[3][30][0]=94;
		input_array[4][30][0]=82;
		input_array[5][30][0]=81;
		input_array[6][30][0]=95;
		input_array[7][30][0]=94;
		input_array[8][30][0]=96;
		input_array[9][30][0]=104;
		input_array[10][30][0]=108;
		input_array[11][30][0]=112;
		input_array[12][30][0]=110;
		input_array[13][30][0]=108;
		input_array[14][30][0]=124;
		input_array[15][30][0]=119;
		input_array[16][30][0]=105;
		input_array[17][30][0]=107;
		input_array[18][30][0]=117;
		input_array[19][30][0]=127;
		input_array[20][30][0]=116;
		input_array[21][30][0]=124;
		input_array[22][30][0]=115;
		input_array[23][30][0]=111;
		input_array[24][30][0]=116;
		input_array[25][30][0]=107;
		input_array[26][30][0]=109;
		input_array[27][30][0]=106;
		input_array[28][30][0]=96;
		input_array[29][30][0]=80;
		input_array[30][30][0]=76;
		input_array[31][30][0]=82;
		input_array[0][31][0]=97;
		input_array[1][31][0]=94;
		input_array[2][31][0]=93;
		input_array[3][31][0]=97;
		input_array[4][31][0]=96;
		input_array[5][31][0]=94;
		input_array[6][31][0]=96;
		input_array[7][31][0]=79;
		input_array[8][31][0]=78;
		input_array[9][31][0]=93;
		input_array[10][31][0]=105;
		input_array[11][31][0]=107;
		input_array[12][31][0]=98;
		input_array[13][31][0]=99;
		input_array[14][31][0]=106;
		input_array[15][31][0]=119;
		input_array[16][31][0]=104;
		input_array[17][31][0]=104;
		input_array[18][31][0]=106;
		input_array[19][31][0]=122;
		input_array[20][31][0]=107;
		input_array[21][31][0]=112;
		input_array[22][31][0]=92;
		input_array[23][31][0]=80;
		input_array[24][31][0]=96;
		input_array[25][31][0]=77;
		input_array[26][31][0]=85;
		input_array[27][31][0]=84;
		input_array[28][31][0]=67;
		input_array[29][31][0]=54;
		input_array[30][31][0]=63;
		input_array[31][31][0]=72;
		input_array[0][0][1]=25;
		input_array[1][0][1]=34;
		input_array[2][0][1]=35;
		input_array[3][0][1]=37;
		input_array[4][0][1]=39;
		input_array[5][0][1]=37;
		input_array[6][0][1]=38;
		input_array[7][0][1]=23;
		input_array[8][0][1]=25;
		input_array[9][0][1]=27;
		input_array[10][0][1]=20;
		input_array[11][0][1]=30;
		input_array[12][0][1]=37;
		input_array[13][0][1]=48;
		input_array[14][0][1]=63;
		input_array[15][0][1]=46;
		input_array[16][0][1]=35;
		input_array[17][0][1]=35;
		input_array[18][0][1]=29;
		input_array[19][0][1]=30;
		input_array[20][0][1]=34;
		input_array[21][0][1]=39;
		input_array[22][0][1]=50;
		input_array[23][0][1]=71;
		input_array[24][0][1]=48;
		input_array[25][0][1]=42;
		input_array[26][0][1]=56;
		input_array[27][0][1]=51;
		input_array[28][0][1]=40;
		input_array[29][0][1]=67;
		input_array[30][0][1]=72;
		input_array[31][0][1]=76;
		input_array[0][1][1]=28;
		input_array[1][1][1]=30;
		input_array[2][1][1]=27;
		input_array[3][1][1]=33;
		input_array[4][1][1]=29;
		input_array[5][1][1]=33;
		input_array[6][1][1]=34;
		input_array[7][1][1]=36;
		input_array[8][1][1]=47;
		input_array[9][1][1]=34;
		input_array[10][1][1]=18;
		input_array[11][1][1]=35;
		input_array[12][1][1]=47;
		input_array[13][1][1]=57;
		input_array[14][1][1]=69;
		input_array[15][1][1]=37;
		input_array[16][1][1]=34;
		input_array[17][1][1]=42;
		input_array[18][1][1]=56;
		input_array[19][1][1]=39;
		input_array[20][1][1]=48;
		input_array[21][1][1]=73;
		input_array[22][1][1]=73;
		input_array[23][1][1]=95;
		input_array[24][1][1]=80;
		input_array[25][1][1]=51;
		input_array[26][1][1]=61;
		input_array[27][1][1]=72;
		input_array[28][1][1]=62;
		input_array[29][1][1]=82;
		input_array[30][1][1]=82;
		input_array[31][1][1]=72;
		input_array[0][2][1]=32;
		input_array[1][2][1]=33;
		input_array[2][2][1]=50;
		input_array[3][2][1]=41;
		input_array[4][2][1]=38;
		input_array[5][2][1]=34;
		input_array[6][2][1]=33;
		input_array[7][2][1]=60;
		input_array[8][2][1]=81;
		input_array[9][2][1]=45;
		input_array[10][2][1]=38;
		input_array[11][2][1]=64;
		input_array[12][2][1]=60;
		input_array[13][2][1]=61;
		input_array[14][2][1]=78;
		input_array[15][2][1]=52;
		input_array[16][2][1]=55;
		input_array[17][2][1]=70;
		input_array[18][2][1]=81;
		input_array[19][2][1]=58;
		input_array[20][2][1]=81;
		input_array[21][2][1]=87;
		input_array[22][2][1]=73;
		input_array[23][2][1]=94;
		input_array[24][2][1]=96;
		input_array[25][2][1]=76;
		input_array[26][2][1]=80;
		input_array[27][2][1]=85;
		input_array[28][2][1]=75;
		input_array[29][2][1]=76;
		input_array[30][2][1]=89;
		input_array[31][2][1]=77;
		input_array[0][3][1]=46;
		input_array[1][3][1]=55;
		input_array[2][3][1]=77;
		input_array[3][3][1]=58;
		input_array[4][3][1]=65;
		input_array[5][3][1]=48;
		input_array[6][3][1]=68;
		input_array[7][3][1]=75;
		input_array[8][3][1]=90;
		input_array[9][3][1]=74;
		input_array[10][3][1]=85;
		input_array[11][3][1]=79;
		input_array[12][3][1]=79;
		input_array[13][3][1]=85;
		input_array[14][3][1]=76;
		input_array[15][3][1]=78;
		input_array[16][3][1]=83;
		input_array[17][3][1]=90;
		input_array[18][3][1]=84;
		input_array[19][3][1]=77;
		input_array[20][3][1]=83;
		input_array[21][3][1]=80;
		input_array[22][3][1]=87;
		input_array[23][3][1]=87;
		input_array[24][3][1]=72;
		input_array[25][3][1]=65;
		input_array[26][3][1]=85;
		input_array[27][3][1]=96;
		input_array[28][3][1]=86;
		input_array[29][3][1]=80;
		input_array[30][3][1]=78;
		input_array[31][3][1]=70;
		input_array[0][4][1]=66;
		input_array[1][4][1]=64;
		input_array[2][4][1]=69;
		input_array[3][4][1]=82;
		input_array[4][4][1]=90;
		input_array[5][4][1]=68;
		input_array[6][4][1]=89;
		input_array[7][4][1]=84;
		input_array[8][4][1]=70;
		input_array[9][4][1]=84;
		input_array[10][4][1]=90;
		input_array[11][4][1]=79;
		input_array[12][4][1]=83;
		input_array[13][4][1]=87;
		input_array[14][4][1]=66;
		input_array[15][4][1]=67;
		input_array[16][4][1]=75;
		input_array[17][4][1]=77;
		input_array[18][4][1]=71;
		input_array[19][4][1]=78;
		input_array[20][4][1]=69;
		input_array[21][4][1]=81;
		input_array[22][4][1]=84;
		input_array[23][4][1]=66;
		input_array[24][4][1]=71;
		input_array[25][4][1]=66;
		input_array[26][4][1]=79;
		input_array[27][4][1]=73;
		input_array[28][4][1]=73;
		input_array[29][4][1]=59;
		input_array[30][4][1]=53;
		input_array[31][4][1]=64;
		input_array[0][5][1]=66;
		input_array[1][5][1]=57;
		input_array[2][5][1]=58;
		input_array[3][5][1]=71;
		input_array[4][5][1]=74;
		input_array[5][5][1]=71;
		input_array[6][5][1]=73;
		input_array[7][5][1]=73;
		input_array[8][5][1]=67;
		input_array[9][5][1]=59;
		input_array[10][5][1]=71;
		input_array[11][5][1]=75;
		input_array[12][5][1]=72;
		input_array[13][5][1]=71;
		input_array[14][5][1]=74;
		input_array[15][5][1]=70;
		input_array[16][5][1]=69;
		input_array[17][5][1]=71;
		input_array[18][5][1]=67;
		input_array[19][5][1]=74;
		input_array[20][5][1]=75;
		input_array[21][5][1]=80;
		input_array[22][5][1]=75;
		input_array[23][5][1]=73;
		input_array[24][5][1]=78;
		input_array[25][5][1]=79;
		input_array[26][5][1]=86;
		input_array[27][5][1]=63;
		input_array[28][5][1]=47;
		input_array[29][5][1]=55;
		input_array[30][5][1]=56;
		input_array[31][5][1]=78;
		input_array[0][6][1]=66;
		input_array[1][6][1]=63;
		input_array[2][6][1]=62;
		input_array[3][6][1]=68;
		input_array[4][6][1]=63;
		input_array[5][6][1]=72;
		input_array[6][6][1]=75;
		input_array[7][6][1]=77;
		input_array[8][6][1]=67;
		input_array[9][6][1]=66;
		input_array[10][6][1]=64;
		input_array[11][6][1]=57;
		input_array[12][6][1]=69;
		input_array[13][6][1]=75;
		input_array[14][6][1]=80;
		input_array[15][6][1]=70;
		input_array[16][6][1]=77;
		input_array[17][6][1]=71;
		input_array[18][6][1]=81;
		input_array[19][6][1]=89;
		input_array[20][6][1]=90;
		input_array[21][6][1]=78;
		input_array[22][6][1]=69;
		input_array[23][6][1]=74;
		input_array[24][6][1]=86;
		input_array[25][6][1]=81;
		input_array[26][6][1]=76;
		input_array[27][6][1]=57;
		input_array[28][6][1]=51;
		input_array[29][6][1]=73;
		input_array[30][6][1]=68;
		input_array[31][6][1]=67;
		input_array[0][7][1]=68;
		input_array[1][7][1]=64;
		input_array[2][7][1]=74;
		input_array[3][7][1]=75;
		input_array[4][7][1]=79;
		input_array[5][7][1]=68;
		input_array[6][7][1]=73;
		input_array[7][7][1]=98;
		input_array[8][7][1]=79;
		input_array[9][7][1]=75;
		input_array[10][7][1]=81;
		input_array[11][7][1]=68;
		input_array[12][7][1]=93;
		input_array[13][7][1]=83;
		input_array[14][7][1]=83;
		input_array[15][7][1]=93;
		input_array[16][7][1]=81;
		input_array[17][7][1]=78;
		input_array[18][7][1]=86;
		input_array[19][7][1]=96;
		input_array[20][7][1]=87;
		input_array[21][7][1]=84;
		input_array[22][7][1]=84;
		input_array[23][7][1]=73;
		input_array[24][7][1]=81;
		input_array[25][7][1]=78;
		input_array[26][7][1]=68;
		input_array[27][7][1]=55;
		input_array[28][7][1]=59;
		input_array[29][7][1]=79;
		input_array[30][7][1]=68;
		input_array[31][7][1]=47;
		input_array[0][8][1]=47;
		input_array[1][8][1]=46;
		input_array[2][8][1]=57;
		input_array[3][8][1]=72;
		input_array[4][8][1]=69;
		input_array[5][8][1]=71;
		input_array[6][8][1]=98;
		input_array[7][8][1]=108;
		input_array[8][8][1]=81;
		input_array[9][8][1]=85;
		input_array[10][8][1]=95;
		input_array[11][8][1]=105;
		input_array[12][8][1]=107;
		input_array[13][8][1]=69;
		input_array[14][8][1]=85;
		input_array[15][8][1]=82;
		input_array[16][8][1]=71;
		input_array[17][8][1]=74;
		input_array[18][8][1]=72;
		input_array[19][8][1]=79;
		input_array[20][8][1]=80;
		input_array[21][8][1]=85;
		input_array[22][8][1]=73;
		input_array[23][8][1]=64;
		input_array[24][8][1]=70;
		input_array[25][8][1]=86;
		input_array[26][8][1]=92;
		input_array[27][8][1]=55;
		input_array[28][8][1]=76;
		input_array[29][8][1]=82;
		input_array[30][8][1]=79;
		input_array[31][8][1]=63;
		input_array[0][9][1]=43;
		input_array[1][9][1]=25;
		input_array[2][9][1]=36;
		input_array[3][9][1]=52;
		input_array[4][9][1]=52;
		input_array[5][9][1]=64;
		input_array[6][9][1]=88;
		input_array[7][9][1]=88;
		input_array[8][9][1]=82;
		input_array[9][9][1]=81;
		input_array[10][9][1]=82;
		input_array[11][9][1]=108;
		input_array[12][9][1]=71;
		input_array[13][9][1]=77;
		input_array[14][9][1]=94;
		input_array[15][9][1]=87;
		input_array[16][9][1]=96;
		input_array[17][9][1]=93;
		input_array[18][9][1]=83;
		input_array[19][9][1]=87;
		input_array[20][9][1]=79;
		input_array[21][9][1]=92;
		input_array[22][9][1]=62;
		input_array[23][9][1]=60;
		input_array[24][9][1]=79;
		input_array[25][9][1]=77;
		input_array[26][9][1]=81;
		input_array[27][9][1]=63;
		input_array[28][9][1]=87;
		input_array[29][9][1]=74;
		input_array[30][9][1]=67;
		input_array[31][9][1]=75;
		input_array[0][10][1]=61;
		input_array[1][10][1]=35;
		input_array[2][10][1]=48;
		input_array[3][10][1]=48;
		input_array[4][10][1]=52;
		input_array[5][10][1]=73;
		input_array[6][10][1]=87;
		input_array[7][10][1]=78;
		input_array[8][10][1]=74;
		input_array[9][10][1]=82;
		input_array[10][10][1]=121;
		input_array[11][10][1]=97;
		input_array[12][10][1]=64;
		input_array[13][10][1]=92;
		input_array[14][10][1]=91;
		input_array[15][10][1]=87;
		input_array[16][10][1]=108;
		input_array[17][10][1]=98;
		input_array[18][10][1]=92;
		input_array[19][10][1]=94;
		input_array[20][10][1]=69;
		input_array[21][10][1]=69;
		input_array[22][10][1]=76;
		input_array[23][10][1]=66;
		input_array[24][10][1]=77;
		input_array[25][10][1]=82;
		input_array[26][10][1]=78;
		input_array[27][10][1]=93;
		input_array[28][10][1]=93;
		input_array[29][10][1]=60;
		input_array[30][10][1]=58;
		input_array[31][10][1]=85;
		input_array[0][11][1]=68;
		input_array[1][11][1]=70;
		input_array[2][11][1]=80;
		input_array[3][11][1]=83;
		input_array[4][11][1]=54;
		input_array[5][11][1]=69;
		input_array[6][11][1]=99;
		input_array[7][11][1]=75;
		input_array[8][11][1]=75;
		input_array[9][11][1]=82;
		input_array[10][11][1]=106;
		input_array[11][11][1]=75;
		input_array[12][11][1]=59;
		input_array[13][11][1]=92;
		input_array[14][11][1]=79;
		input_array[15][11][1]=78;
		input_array[16][11][1]=98;
		input_array[17][11][1]=84;
		input_array[18][11][1]=94;
		input_array[19][11][1]=94;
		input_array[20][11][1]=70;
		input_array[21][11][1]=72;
		input_array[22][11][1]=89;
		input_array[23][11][1]=86;
		input_array[24][11][1]=90;
		input_array[25][11][1]=103;
		input_array[26][11][1]=105;
		input_array[27][11][1]=103;
		input_array[28][11][1]=73;
		input_array[29][11][1]=64;
		input_array[30][11][1]=67;
		input_array[31][11][1]=75;
		input_array[0][12][1]=74;
		input_array[1][12][1]=84;
		input_array[2][12][1]=90;
		input_array[3][12][1]=106;
		input_array[4][12][1]=84;
		input_array[5][12][1]=65;
		input_array[6][12][1]=58;
		input_array[7][12][1]=56;
		input_array[8][12][1]=62;
		input_array[9][12][1]=86;
		input_array[10][12][1]=79;
		input_array[11][12][1]=55;
		input_array[12][12][1]=51;
		input_array[13][12][1]=77;
		input_array[14][12][1]=78;
		input_array[15][12][1]=76;
		input_array[16][12][1]=82;
		input_array[17][12][1]=76;
		input_array[18][12][1]=77;
		input_array[19][12][1]=87;
		input_array[20][12][1]=89;
		input_array[21][12][1]=90;
		input_array[22][12][1]=86;
		input_array[23][12][1]=84;
		input_array[24][12][1]=82;
		input_array[25][12][1]=90;
		input_array[26][12][1]=86;
		input_array[27][12][1]=79;
		input_array[28][12][1]=71;
		input_array[29][12][1]=74;
		input_array[30][12][1]=74;
		input_array[31][12][1]=80;
		input_array[0][13][1]=98;
		input_array[1][13][1]=96;
		input_array[2][13][1]=112;
		input_array[3][13][1]=113;
		input_array[4][13][1]=104;
		input_array[5][13][1]=105;
		input_array[6][13][1]=40;
		input_array[7][13][1]=38;
		input_array[8][13][1]=51;
		input_array[9][13][1]=61;
		input_array[10][13][1]=78;
		input_array[11][13][1]=70;
		input_array[12][13][1]=48;
		input_array[13][13][1]=55;
		input_array[14][13][1]=72;
		input_array[15][13][1]=83;
		input_array[16][13][1]=100;
		input_array[17][13][1]=111;
		input_array[18][13][1]=126;
		input_array[19][13][1]=138;
		input_array[20][13][1]=129;
		input_array[21][13][1]=93;
		input_array[22][13][1]=94;
		input_array[23][13][1]=87;
		input_array[24][13][1]=78;
		input_array[25][13][1]=83;
		input_array[26][13][1]=86;
		input_array[27][13][1]=79;
		input_array[28][13][1]=79;
		input_array[29][13][1]=80;
		input_array[30][13][1]=75;
		input_array[31][13][1]=73;
		input_array[0][14][1]=97;
		input_array[1][14][1]=102;
		input_array[2][14][1]=115;
		input_array[3][14][1]=104;
		input_array[4][14][1]=107;
		input_array[5][14][1]=112;
		input_array[6][14][1]=38;
		input_array[7][14][1]=40;
		input_array[8][14][1]=51;
		input_array[9][14][1]=59;
		input_array[10][14][1]=109;
		input_array[11][14][1]=130;
		input_array[12][14][1]=105;
		input_array[13][14][1]=112;
		input_array[14][14][1]=127;
		input_array[15][14][1]=130;
		input_array[16][14][1]=108;
		input_array[17][14][1]=166;
		input_array[18][14][1]=192;
		input_array[19][14][1]=191;
		input_array[20][14][1]=172;
		input_array[21][14][1]=109;
		input_array[22][14][1]=93;
		input_array[23][14][1]=90;
		input_array[24][14][1]=98;
		input_array[25][14][1]=96;
		input_array[26][14][1]=93;
		input_array[27][14][1]=98;
		input_array[28][14][1]=83;
		input_array[29][14][1]=85;
		input_array[30][14][1]=71;
		input_array[31][14][1]=66;
		input_array[0][15][1]=68;
		input_array[1][15][1]=79;
		input_array[2][15][1]=89;
		input_array[3][15][1]=96;
		input_array[4][15][1]=96;
		input_array[5][15][1]=100;
		input_array[6][15][1]=51;
		input_array[7][15][1]=42;
		input_array[8][15][1]=72;
		input_array[9][15][1]=74;
		input_array[10][15][1]=143;
		input_array[11][15][1]=150;
		input_array[12][15][1]=135;
		input_array[13][15][1]=142;
		input_array[14][15][1]=151;
		input_array[15][15][1]=153;
		input_array[16][15][1]=121;
		input_array[17][15][1]=152;
		input_array[18][15][1]=181;
		input_array[19][15][1]=206;
		input_array[20][15][1]=187;
		input_array[21][15][1]=138;
		input_array[22][15][1]=117;
		input_array[23][15][1]=106;
		input_array[24][15][1]=112;
		input_array[25][15][1]=113;
		input_array[26][15][1]=108;
		input_array[27][15][1]=112;
		input_array[28][15][1]=91;
		input_array[29][15][1]=99;
		input_array[30][15][1]=81;
		input_array[31][15][1]=92;
		input_array[0][16][1]=59;
		input_array[1][16][1]=68;
		input_array[2][16][1]=75;
		input_array[3][16][1]=96;
		input_array[4][16][1]=94;
		input_array[5][16][1]=92;
		input_array[6][16][1]=80;
		input_array[7][16][1]=36;
		input_array[8][16][1]=76;
		input_array[9][16][1]=100;
		input_array[10][16][1]=164;
		input_array[11][16][1]=165;
		input_array[12][16][1]=155;
		input_array[13][16][1]=162;
		input_array[14][16][1]=172;
		input_array[15][16][1]=175;
		input_array[16][16][1]=144;
		input_array[17][16][1]=138;
		input_array[18][16][1]=160;
		input_array[19][16][1]=183;
		input_array[20][16][1]=191;
		input_array[21][16][1]=148;
		input_array[22][16][1]=130;
		input_array[23][16][1]=107;
		input_array[24][16][1]=109;
		input_array[25][16][1]=117;
		input_array[26][16][1]=117;
		input_array[27][16][1]=112;
		input_array[28][16][1]=100;
		input_array[29][16][1]=104;
		input_array[30][16][1]=91;
		input_array[31][16][1]=95;
		input_array[0][17][1]=62;
		input_array[1][17][1]=60;
		input_array[2][17][1]=72;
		input_array[3][17][1]=90;
		input_array[4][17][1]=98;
		input_array[5][17][1]=93;
		input_array[6][17][1]=74;
		input_array[7][17][1]=19;
		input_array[8][17][1]=64;
		input_array[9][17][1]=130;
		input_array[10][17][1]=171;
		input_array[11][17][1]=181;
		input_array[12][17][1]=182;
		input_array[13][17][1]=178;
		input_array[14][17][1]=175;
		input_array[15][17][1]=178;
		input_array[16][17][1]=164;
		input_array[17][17][1]=142;
		input_array[18][17][1]=139;
		input_array[19][17][1]=116;
		input_array[20][17][1]=152;
		input_array[21][17][1]=127;
		input_array[22][17][1]=102;
		input_array[23][17][1]=102;
		input_array[24][17][1]=116;
		input_array[25][17][1]=117;
		input_array[26][17][1]=124;
		input_array[27][17][1]=121;
		input_array[28][17][1]=104;
		input_array[29][17][1]=105;
		input_array[30][17][1]=109;
		input_array[31][17][1]=97;
		input_array[0][18][1]=82;
		input_array[1][18][1]=87;
		input_array[2][18][1]=94;
		input_array[3][18][1]=104;
		input_array[4][18][1]=101;
		input_array[5][18][1]=96;
		input_array[6][18][1]=82;
		input_array[7][18][1]=46;
		input_array[8][18][1]=74;
		input_array[9][18][1]=152;
		input_array[10][18][1]=178;
		input_array[11][18][1]=192;
		input_array[12][18][1]=194;
		input_array[13][18][1]=192;
		input_array[14][18][1]=177;
		input_array[15][18][1]=189;
		input_array[16][18][1]=188;
		input_array[17][18][1]=143;
		input_array[18][18][1]=121;
		input_array[19][18][1]=80;
		input_array[20][18][1]=94;
		input_array[21][18][1]=79;
		input_array[22][18][1]=74;
		input_array[23][18][1]=115;
		input_array[24][18][1]=124;
		input_array[25][18][1]=114;
		input_array[26][18][1]=122;
		input_array[27][18][1]=120;
		input_array[28][18][1]=110;
		input_array[29][18][1]=106;
		input_array[30][18][1]=112;
		input_array[31][18][1]=94;
		input_array[0][19][1]=84;
		input_array[1][19][1]=96;
		input_array[2][19][1]=100;
		input_array[3][19][1]=111;
		input_array[4][19][1]=98;
		input_array[5][19][1]=91;
		input_array[6][19][1]=95;
		input_array[7][19][1]=94;
		input_array[8][19][1]=99;
		input_array[9][19][1]=157;
		input_array[10][19][1]=182;
		input_array[11][19][1]=190;
		input_array[12][19][1]=194;
		input_array[13][19][1]=198;
		input_array[14][19][1]=189;
		input_array[15][19][1]=196;
		input_array[16][19][1]=194;
		input_array[17][19][1]=145;
		input_array[18][19][1]=81;
		input_array[19][19][1]=70;
		input_array[20][19][1]=77;
		input_array[21][19][1]=70;
		input_array[22][19][1]=73;
		input_array[23][19][1]=117;
		input_array[24][19][1]=125;
		input_array[25][19][1]=116;
		input_array[26][19][1]=113;
		input_array[27][19][1]=103;
		input_array[28][19][1]=106;
		input_array[29][19][1]=100;
		input_array[30][19][1]=99;
		input_array[31][19][1]=87;
		input_array[0][20][1]=79;
		input_array[1][20][1]=85;
		input_array[2][20][1]=98;
		input_array[3][20][1]=95;
		input_array[4][20][1]=91;
		input_array[5][20][1]=100;
		input_array[6][20][1]=102;
		input_array[7][20][1]=83;
		input_array[8][20][1]=88;
		input_array[9][20][1]=145;
		input_array[10][20][1]=179;
		input_array[11][20][1]=183;
		input_array[12][20][1]=194;
		input_array[13][20][1]=200;
		input_array[14][20][1]=186;
		input_array[15][20][1]=193;
		input_array[16][20][1]=184;
		input_array[17][20][1]=152;
		input_array[18][20][1]=57;
		input_array[19][20][1]=56;
		input_array[20][20][1]=59;
		input_array[21][20][1]=63;
		input_array[22][20][1]=71;
		input_array[23][20][1]=107;
		input_array[24][20][1]=111;
		input_array[25][20][1]=117;
		input_array[26][20][1]=105;
		input_array[27][20][1]=84;
		input_array[28][20][1]=84;
		input_array[29][20][1]=83;
		input_array[30][20][1]=84;
		input_array[31][20][1]=91;
		input_array[0][21][1]=62;
		input_array[1][21][1]=84;
		input_array[2][21][1]=87;
		input_array[3][21][1]=85;
		input_array[4][21][1]=104;
		input_array[5][21][1]=90;
		input_array[6][21][1]=86;
		input_array[7][21][1]=77;
		input_array[8][21][1]=82;
		input_array[9][21][1]=109;
		input_array[10][21][1]=146;
		input_array[11][21][1]=149;
		input_array[12][21][1]=181;
		input_array[13][21][1]=193;
		input_array[14][21][1]=175;
		input_array[15][21][1]=180;
		input_array[16][21][1]=174;
		input_array[17][21][1]=155;
		input_array[18][21][1]=40;
		input_array[19][21][1]=13;
		input_array[20][21][1]=34;
		input_array[21][21][1]=47;
		input_array[22][21][1]=65;
		input_array[23][21][1]=96;
		input_array[24][21][1]=92;
		input_array[25][21][1]=98;
		input_array[26][21][1]=89;
		input_array[27][21][1]=75;
		input_array[28][21][1]=74;
		input_array[29][21][1]=74;
		input_array[30][21][1]=75;
		input_array[31][21][1]=74;
		input_array[0][22][1]=36;
		input_array[1][22][1]=67;
		input_array[2][22][1]=61;
		input_array[3][22][1]=90;
		input_array[4][22][1]=94;
		input_array[5][22][1]=78;
		input_array[6][22][1]=74;
		input_array[7][22][1]=76;
		input_array[8][22][1]=78;
		input_array[9][22][1]=73;
		input_array[10][22][1]=111;
		input_array[11][22][1]=82;
		input_array[12][22][1]=100;
		input_array[13][22][1]=115;
		input_array[14][22][1]=78;
		input_array[15][22][1]=78;
		input_array[16][22][1]=153;
		input_array[17][22][1]=152;
		input_array[18][22][1]=56;
		input_array[19][22][1]=26;
		input_array[20][22][1]=18;
		input_array[21][22][1]=28;
		input_array[22][22][1]=52;
		input_array[23][22][1]=84;
		input_array[24][22][1]=77;
		input_array[25][22][1]=71;
		input_array[26][22][1]=77;
		input_array[27][22][1]=70;
		input_array[28][22][1]=73;
		input_array[29][22][1]=71;
		input_array[30][22][1]=59;
		input_array[31][22][1]=72;
		input_array[0][23][1]=35;
		input_array[1][23][1]=52;
		input_array[2][23][1]=62;
		input_array[3][23][1]=78;
		input_array[4][23][1]=82;
		input_array[5][23][1]=78;
		input_array[6][23][1]=65;
		input_array[7][23][1]=67;
		input_array[8][23][1]=65;
		input_array[9][23][1]=74;
		input_array[10][23][1]=93;
		input_array[11][23][1]=37;
		input_array[12][23][1]=46;
		input_array[13][23][1]=38;
		input_array[14][23][1]=38;
		input_array[15][23][1]=46;
		input_array[16][23][1]=116;
		input_array[17][23][1]=126;
		input_array[18][23][1]=67;
		input_array[19][23][1]=50;
		input_array[20][23][1]=19;
		input_array[21][23][1]=32;
		input_array[22][23][1]=31;
		input_array[23][23][1]=80;
		input_array[24][23][1]=75;
		input_array[25][23][1]=67;
		input_array[26][23][1]=60;
		input_array[27][23][1]=58;
		input_array[28][23][1]=56;
		input_array[29][23][1]=70;
		input_array[30][23][1]=57;
		input_array[31][23][1]=66;
		input_array[0][24][1]=54;
		input_array[1][24][1]=68;
		input_array[2][24][1]=73;
		input_array[3][24][1]=64;
		input_array[4][24][1]=73;
		input_array[5][24][1]=67;
		input_array[6][24][1]=61;
		input_array[7][24][1]=66;
		input_array[8][24][1]=72;
		input_array[9][24][1]=71;
		input_array[10][24][1]=75;
		input_array[11][24][1]=33;
		input_array[12][24][1]=59;
		input_array[13][24][1]=80;
		input_array[14][24][1]=75;
		input_array[15][24][1]=62;
		input_array[16][24][1]=88;
		input_array[17][24][1]=109;
		input_array[18][24][1]=66;
		input_array[19][24][1]=60;
		input_array[20][24][1]=41;
		input_array[21][24][1]=50;
		input_array[22][24][1]=34;
		input_array[23][24][1]=49;
		input_array[24][24][1]=87;
		input_array[25][24][1]=74;
		input_array[26][24][1]=64;
		input_array[27][24][1]=62;
		input_array[28][24][1]=51;
		input_array[29][24][1]=88;
		input_array[30][24][1]=78;
		input_array[31][24][1]=69;
		input_array[0][25][1]=44;
		input_array[1][25][1]=52;
		input_array[2][25][1]=75;
		input_array[3][25][1]=73;
		input_array[4][25][1]=66;
		input_array[5][25][1]=76;
		input_array[6][25][1]=71;
		input_array[7][25][1]=74;
		input_array[8][25][1]=80;
		input_array[9][25][1]=76;
		input_array[10][25][1]=67;
		input_array[11][25][1]=42;
		input_array[12][25][1]=78;
		input_array[13][25][1]=82;
		input_array[14][25][1]=79;
		input_array[15][25][1]=78;
		input_array[16][25][1]=92;
		input_array[17][25][1]=97;
		input_array[18][25][1]=100;
		input_array[19][25][1]=76;
		input_array[20][25][1]=49;
		input_array[21][25][1]=38;
		input_array[22][25][1]=70;
		input_array[23][25][1]=41;
		input_array[24][25][1]=83;
		input_array[25][25][1]=74;
		input_array[26][25][1]=50;
		input_array[27][25][1]=50;
		input_array[28][25][1]=60;
		input_array[29][25][1]=98;
		input_array[30][25][1]=77;
		input_array[31][25][1]=79;
		input_array[0][26][1]=55;
		input_array[1][26][1]=51;
		input_array[2][26][1]=70;
		input_array[3][26][1]=75;
		input_array[4][26][1]=71;
		input_array[5][26][1]=79;
		input_array[6][26][1]=76;
		input_array[7][26][1]=81;
		input_array[8][26][1]=86;
		input_array[9][26][1]=80;
		input_array[10][26][1]=65;
		input_array[11][26][1]=46;
		input_array[12][26][1]=93;
		input_array[13][26][1]=80;
		input_array[14][26][1]=88;
		input_array[15][26][1]=67;
		input_array[16][26][1]=82;
		input_array[17][26][1]=91;
		input_array[18][26][1]=107;
		input_array[19][26][1]=84;
		input_array[20][26][1]=70;
		input_array[21][26][1]=48;
		input_array[22][26][1]=80;
		input_array[23][26][1]=63;
		input_array[24][26][1]=69;
		input_array[25][26][1]=66;
		input_array[26][26][1]=51;
		input_array[27][26][1]=66;
		input_array[28][26][1]=80;
		input_array[29][26][1]=83;
		input_array[30][26][1]=57;
		input_array[31][26][1]=59;
		input_array[0][27][1]=64;
		input_array[1][27][1]=65;
		input_array[2][27][1]=64;
		input_array[3][27][1]=68;
		input_array[4][27][1]=75;
		input_array[5][27][1]=79;
		input_array[6][27][1]=81;
		input_array[7][27][1]=84;
		input_array[8][27][1]=101;
		input_array[9][27][1]=87;
		input_array[10][27][1]=69;
		input_array[11][27][1]=53;
		input_array[12][27][1]=87;
		input_array[13][27][1]=83;
		input_array[14][27][1]=81;
		input_array[15][27][1]=58;
		input_array[16][27][1]=59;
		input_array[17][27][1]=86;
		input_array[18][27][1]=82;
		input_array[19][27][1]=83;
		input_array[20][27][1]=83;
		input_array[21][27][1]=85;
		input_array[22][27][1]=66;
		input_array[23][27][1]=78;
		input_array[24][27][1]=80;
		input_array[25][27][1]=76;
		input_array[26][27][1]=91;
		input_array[27][27][1]=90;
		input_array[28][27][1]=80;
		input_array[29][27][1]=72;
		input_array[30][27][1]=72;
		input_array[31][27][1]=68;
		input_array[0][28][1]=67;
		input_array[1][28][1]=77;
		input_array[2][28][1]=74;
		input_array[3][28][1]=74;
		input_array[4][28][1]=78;
		input_array[5][28][1]=76;
		input_array[6][28][1]=75;
		input_array[7][28][1]=78;
		input_array[8][28][1]=88;
		input_array[9][28][1]=73;
		input_array[10][28][1]=69;
		input_array[11][28][1]=61;
		input_array[12][28][1]=82;
		input_array[13][28][1]=73;
		input_array[14][28][1]=58;
		input_array[15][28][1]=62;
		input_array[16][28][1]=80;
		input_array[17][28][1]=92;
		input_array[18][28][1]=76;
		input_array[19][28][1]=82;
		input_array[20][28][1]=89;
		input_array[21][28][1]=94;
		input_array[22][28][1]=80;
		input_array[23][28][1]=84;
		input_array[24][28][1]=102;
		input_array[25][28][1]=88;
		input_array[26][28][1]=93;
		input_array[27][28][1]=80;
		input_array[28][28][1]=70;
		input_array[29][28][1]=80;
		input_array[30][28][1]=81;
		input_array[31][28][1]=80;
		input_array[0][29][1]=73;
		input_array[1][29][1]=77;
		input_array[2][29][1]=74;
		input_array[3][29][1]=82;
		input_array[4][29][1]=70;
		input_array[5][29][1]=73;
		input_array[6][29][1]=80;
		input_array[7][29][1]=91;
		input_array[8][29][1]=98;
		input_array[9][29][1]=90;
		input_array[10][29][1]=75;
		input_array[11][29][1]=91;
		input_array[12][29][1]=91;
		input_array[13][29][1]=93;
		input_array[14][29][1]=94;
		input_array[15][29][1]=92;
		input_array[16][29][1]=92;
		input_array[17][29][1]=89;
		input_array[18][29][1]=88;
		input_array[19][29][1]=98;
		input_array[20][29][1]=99;
		input_array[21][29][1]=100;
		input_array[22][29][1]=101;
		input_array[23][29][1]=99;
		input_array[24][29][1]=106;
		input_array[25][29][1]=95;
		input_array[26][29][1]=94;
		input_array[27][29][1]=90;
		input_array[28][29][1]=90;
		input_array[29][29][1]=93;
		input_array[30][29][1]=84;
		input_array[31][29][1]=75;
		input_array[0][30][1]=72;
		input_array[1][30][1]=74;
		input_array[2][30][1]=77;
		input_array[3][30][1]=82;
		input_array[4][30][1]=72;
		input_array[5][30][1]=71;
		input_array[6][30][1]=85;
		input_array[7][30][1]=87;
		input_array[8][30][1]=89;
		input_array[9][30][1]=91;
		input_array[10][30][1]=88;
		input_array[11][30][1]=92;
		input_array[12][30][1]=98;
		input_array[13][30][1]=92;
		input_array[14][30][1]=105;
		input_array[15][30][1]=98;
		input_array[16][30][1]=89;
		input_array[17][30][1]=85;
		input_array[18][30][1]=91;
		input_array[19][30][1]=104;
		input_array[20][30][1]=94;
		input_array[21][30][1]=107;
		input_array[22][30][1]=101;
		input_array[23][30][1]=92;
		input_array[24][30][1]=98;
		input_array[25][30][1]=97;
		input_array[26][30][1]=100;
		input_array[27][30][1]=96;
		input_array[28][30][1]=87;
		input_array[29][30][1]=74;
		input_array[30][30][1]=70;
		input_array[31][30][1]=76;
		input_array[0][31][1]=78;
		input_array[1][31][1]=75;
		input_array[2][31][1]=75;
		input_array[3][31][1]=85;
		input_array[4][31][1]=86;
		input_array[5][31][1]=84;
		input_array[6][31][1]=86;
		input_array[7][31][1]=71;
		input_array[8][31][1]=69;
		input_array[9][31][1]=78;
		input_array[10][31][1]=84;
		input_array[11][31][1]=86;
		input_array[12][31][1]=85;
		input_array[13][31][1]=83;
		input_array[14][31][1]=87;
		input_array[15][31][1]=98;
		input_array[16][31][1]=88;
		input_array[17][31][1]=85;
		input_array[18][31][1]=85;
		input_array[19][31][1]=99;
		input_array[20][31][1]=85;
		input_array[21][31][1]=96;
		input_array[22][31][1]=81;
		input_array[23][31][1]=62;
		input_array[24][31][1]=78;
		input_array[25][31][1]=67;
		input_array[26][31][1]=76;
		input_array[27][31][1]=75;
		input_array[28][31][1]=57;
		input_array[29][31][1]=47;
		input_array[30][31][1]=56;
		input_array[31][31][1]=65;
		input_array[0][0][2]=10;
		input_array[1][0][2]=19;
		input_array[2][0][2]=20;
		input_array[3][0][2]=23;
		input_array[4][0][2]=25;
		input_array[5][0][2]=22;
		input_array[6][0][2]=23;
		input_array[7][0][2]=9;
		input_array[8][0][2]=15;
		input_array[9][0][2]=19;
		input_array[10][0][2]=10;
		input_array[11][0][2]=17;
		input_array[12][0][2]=23;
		input_array[13][0][2]=34;
		input_array[14][0][2]=50;
		input_array[15][0][2]=32;
		input_array[16][0][2]=25;
		input_array[17][0][2]=25;
		input_array[18][0][2]=20;
		input_array[19][0][2]=20;
		input_array[20][0][2]=23;
		input_array[21][0][2]=25;
		input_array[22][0][2]=33;
		input_array[23][0][2]=50;
		input_array[24][0][2]=27;
		input_array[25][0][2]=24;
		input_array[26][0][2]=41;
		input_array[27][0][2]=40;
		input_array[28][0][2]=25;
		input_array[29][0][2]=39;
		input_array[30][0][2]=43;
		input_array[31][0][2]=47;
		input_array[0][1][2]=13;
		input_array[1][1][2]=14;
		input_array[2][1][2]=12;
		input_array[3][1][2]=18;
		input_array[4][1][2]=14;
		input_array[5][1][2]=17;
		input_array[6][1][2]=18;
		input_array[7][1][2]=19;
		input_array[8][1][2]=30;
		input_array[9][1][2]=19;
		input_array[10][1][2]=4;
		input_array[11][1][2]=19;
		input_array[12][1][2]=32;
		input_array[13][1][2]=42;
		input_array[14][1][2]=55;
		input_array[15][1][2]=25;
		input_array[16][1][2]=18;
		input_array[17][1][2]=25;
		input_array[18][1][2]=40;
		input_array[19][1][2]=23;
		input_array[20][1][2]=31;
		input_array[21][1][2]=53;
		input_array[22][1][2]=52;
		input_array[23][1][2]=70;
		input_array[24][1][2]=58;
		input_array[25][1][2]=32;
		input_array[26][1][2]=42;
		input_array[27][1][2]=52;
		input_array[28][1][2]=40;
		input_array[29][1][2]=55;
		input_array[30][1][2]=56;
		input_array[31][1][2]=45;
		input_array[0][2][2]=15;
		input_array[1][2][2]=17;
		input_array[2][2][2]=33;
		input_array[3][2][2]=23;
		input_array[4][2][2]=21;
		input_array[5][2][2]=17;
		input_array[6][2][2]=17;
		input_array[7][2][2]=40;
		input_array[8][2][2]=59;
		input_array[9][2][2]=24;
		input_array[10][2][2]=19;
		input_array[11][2][2]=43;
		input_array[12][2][2]=45;
		input_array[13][2][2]=46;
		input_array[14][2][2]=63;
		input_array[15][2][2]=38;
		input_array[16][2][2]=34;
		input_array[17][2][2]=49;
		input_array[18][2][2]=59;
		input_array[19][2][2]=36;
		input_array[20][2][2]=56;
		input_array[21][2][2]=61;
		input_array[22][2][2]=46;
		input_array[23][2][2]=65;
		input_array[24][2][2]=73;
		input_array[25][2][2]=57;
		input_array[26][2][2]=57;
		input_array[27][2][2]=56;
		input_array[28][2][2]=47;
		input_array[29][2][2]=52;
		input_array[30][2][2]=66;
		input_array[31][2][2]=54;
		input_array[0][3][2]=28;
		input_array[1][3][2]=36;
		input_array[2][3][2]=58;
		input_array[3][3][2]=39;
		input_array[4][3][2]=46;
		input_array[5][3][2]=30;
		input_array[6][3][2]=51;
		input_array[7][3][2]=54;
		input_array[8][3][2]=64;
		input_array[9][3][2]=48;
		input_array[10][3][2]=59;
		input_array[11][3][2]=55;
		input_array[12][3][2]=61;
		input_array[13][3][2]=68;
		input_array[14][3][2]=59;
		input_array[15][3][2]=60;
		input_array[16][3][2]=58;
		input_array[17][3][2]=64;
		input_array[18][3][2]=58;
		input_array[19][3][2]=51;
		input_array[20][3][2]=54;
		input_array[21][3][2]=50;
		input_array[22][3][2]=56;
		input_array[23][3][2]=56;
		input_array[24][3][2]=48;
		input_array[25][3][2]=45;
		input_array[26][3][2]=58;
		input_array[27][3][2]=61;
		input_array[28][3][2]=53;
		input_array[29][3][2]=59;
		input_array[30][3][2]=57;
		input_array[31][3][2]=49;
		input_array[0][4][2]=47;
		input_array[1][4][2]=45;
		input_array[2][4][2]=50;
		input_array[3][4][2]=61;
		input_array[4][4][2]=70;
		input_array[5][4][2]=49;
		input_array[6][4][2]=72;
		input_array[7][4][2]=62;
		input_array[8][4][2]=42;
		input_array[9][4][2]=55;
		input_array[10][4][2]=61;
		input_array[11][4][2]=53;
		input_array[12][4][2]=62;
		input_array[13][4][2]=67;
		input_array[14][4][2]=45;
		input_array[15][4][2]=45;
		input_array[16][4][2]=48;
		input_array[17][4][2]=49;
		input_array[18][4][2]=42;
		input_array[19][4][2]=49;
		input_array[20][4][2]=38;
		input_array[21][4][2]=48;
		input_array[22][4][2]=53;
		input_array[23][4][2]=36;
		input_array[24][4][2]=47;
		input_array[25][4][2]=45;
		input_array[26][4][2]=51;
		input_array[27][4][2]=39;
		input_array[28][4][2]=40;
		input_array[29][4][2]=37;
		input_array[30][4][2]=32;
		input_array[31][4][2]=43;
		input_array[0][5][2]=45;
		input_array[1][5][2]=37;
		input_array[2][5][2]=38;
		input_array[3][5][2]=48;
		input_array[4][5][2]=51;
		input_array[5][5][2]=51;
		input_array[6][5][2]=54;
		input_array[7][5][2]=51;
		input_array[8][5][2]=39;
		input_array[9][5][2]=30;
		input_array[10][5][2]=43;
		input_array[11][5][2]=49;
		input_array[12][5][2]=47;
		input_array[13][5][2]=46;
		input_array[14][5][2]=49;
		input_array[15][5][2]=44;
		input_array[16][5][2]=41;
		input_array[17][5][2]=43;
		input_array[18][5][2]=39;
		input_array[19][5][2]=46;
		input_array[20][5][2]=43;
		input_array[21][5][2]=48;
		input_array[22][5][2]=46;
		input_array[23][5][2]=46;
		input_array[24][5][2]=54;
		input_array[25][5][2]=55;
		input_array[26][5][2]=61;
		input_array[27][5][2]=35;
		input_array[28][5][2]=20;
		input_array[29][5][2]=35;
		input_array[30][5][2]=35;
		input_array[31][5][2]=58;
		input_array[0][6][2]=44;
		input_array[1][6][2]=41;
		input_array[2][6][2]=40;
		input_array[3][6][2]=43;
		input_array[4][6][2]=39;
		input_array[5][6][2]=50;
		input_array[6][6][2]=55;
		input_array[7][6][2]=56;
		input_array[8][6][2]=42;
		input_array[9][6][2]=38;
		input_array[10][6][2]=37;
		input_array[11][6][2]=32;
		input_array[12][6][2]=41;
		input_array[13][6][2]=47;
		input_array[14][6][2]=52;
		input_array[15][6][2]=42;
		input_array[16][6][2]=50;
		input_array[17][6][2]=45;
		input_array[18][6][2]=55;
		input_array[19][6][2]=63;
		input_array[20][6][2]=60;
		input_array[21][6][2]=48;
		input_array[22][6][2]=43;
		input_array[23][6][2]=50;
		input_array[24][6][2]=62;
		input_array[25][6][2]=57;
		input_array[26][6][2]=54;
		input_array[27][6][2]=37;
		input_array[28][6][2]=32;
		input_array[29][6][2]=53;
		input_array[30][6][2]=49;
		input_array[31][6][2]=48;
		input_array[0][7][2]=46;
		input_array[1][7][2]=43;
		input_array[2][7][2]=52;
		input_array[3][7][2]=50;
		input_array[4][7][2]=54;
		input_array[5][7][2]=47;
		input_array[6][7][2]=54;
		input_array[7][7][2]=78;
		input_array[8][7][2]=55;
		input_array[9][7][2]=49;
		input_array[10][7][2]=56;
		input_array[11][7][2]=44;
		input_array[12][7][2]=62;
		input_array[13][7][2]=52;
		input_array[14][7][2]=52;
		input_array[15][7][2]=63;
		input_array[16][7][2]=57;
		input_array[17][7][2]=55;
		input_array[18][7][2]=62;
		input_array[19][7][2]=72;
		input_array[20][7][2]=60;
		input_array[21][7][2]=57;
		input_array[22][7][2]=60;
		input_array[23][7][2]=53;
		input_array[24][7][2]=59;
		input_array[25][7][2]=53;
		input_array[26][7][2]=48;
		input_array[27][7][2]=40;
		input_array[28][7][2]=45;
		input_array[29][7][2]=59;
		input_array[30][7][2]=47;
		input_array[31][7][2]=26;
		input_array[0][8][2]=31;
		input_array[1][8][2]=30;
		input_array[2][8][2]=41;
		input_array[3][8][2]=52;
		input_array[4][8][2]=51;
		input_array[5][8][2]=55;
		input_array[6][8][2]=72;
		input_array[7][8][2]=79;
		input_array[8][8][2]=55;
		input_array[9][8][2]=55;
		input_array[10][8][2]=64;
		input_array[11][8][2]=76;
		input_array[12][8][2]=75;
		input_array[13][8][2]=36;
		input_array[14][8][2]=50;
		input_array[15][8][2]=46;
		input_array[16][8][2]=42;
		input_array[17][8][2]=50;
		input_array[18][8][2]=51;
		input_array[19][8][2]=55;
		input_array[20][8][2]=58;
		input_array[21][8][2]=60;
		input_array[22][8][2]=47;
		input_array[23][8][2]=47;
		input_array[24][8][2]=52;
		input_array[25][8][2]=62;
		input_array[26][8][2]=70;
		input_array[27][8][2]=36;
		input_array[28][8][2]=57;
		input_array[29][8][2]=59;
		input_array[30][8][2]=56;
		input_array[31][8][2]=39;
		input_array[0][9][2]=29;
		input_array[1][9][2]=11;
		input_array[2][9][2]=22;
		input_array[3][9][2]=35;
		input_array[4][9][2]=39;
		input_array[5][9][2]=50;
		input_array[6][9][2]=58;
		input_array[7][9][2]=54;
		input_array[8][9][2]=54;
		input_array[9][9][2]=50;
		input_array[10][9][2]=48;
		input_array[11][9][2]=76;
		input_array[12][9][2]=42;
		input_array[13][9][2]=46;
		input_array[14][9][2]=59;
		input_array[15][9][2]=50;
		input_array[16][9][2]=64;
		input_array[17][9][2]=69;
		input_array[18][9][2]=62;
		input_array[19][9][2]=62;
		input_array[20][9][2]=59;
		input_array[21][9][2]=68;
		input_array[22][9][2]=34;
		input_array[23][9][2]=43;
		input_array[24][9][2]=63;
		input_array[25][9][2]=53;
		input_array[26][9][2]=57;
		input_array[27][9][2]=39;
		input_array[28][9][2]=63;
		input_array[29][9][2]=51;
		input_array[30][9][2]=43;
		input_array[31][9][2]=51;
		input_array[0][10][2]=42;
		input_array[1][10][2]=17;
		input_array[2][10][2]=29;
		input_array[3][10][2]=29;
		input_array[4][10][2]=37;
		input_array[5][10][2]=56;
		input_array[6][10][2]=58;
		input_array[7][10][2]=48;
		input_array[8][10][2]=50;
		input_array[9][10][2]=54;
		input_array[10][10][2]=90;
		input_array[11][10][2]=67;
		input_array[12][10][2]=41;
		input_array[13][10][2]=67;
		input_array[14][10][2]=62;
		input_array[15][10][2]=55;
		input_array[16][10][2]=75;
		input_array[17][10][2]=73;
		input_array[18][10][2]=70;
		input_array[19][10][2]=67;
		input_array[20][10][2]=47;
		input_array[21][10][2]=44;
		input_array[22][10][2]=48;
		input_array[23][10][2]=47;
		input_array[24][10][2]=58;
		input_array[25][10][2]=58;
		input_array[26][10][2]=54;
		input_array[27][10][2]=68;
		input_array[28][10][2]=69;
		input_array[29][10][2]=39;
		input_array[30][10][2]=37;
		input_array[31][10][2]=64;
		input_array[0][11][2]=45;
		input_array[1][11][2]=47;
		input_array[2][11][2]=57;
		input_array[3][11][2]=61;
		input_array[4][11][2]=36;
		input_array[5][11][2]=49;
		input_array[6][11][2]=71;
		input_array[7][11][2]=50;
		input_array[8][11][2]=56;
		input_array[9][11][2]=57;
		input_array[10][11][2]=77;
		input_array[11][11][2]=47;
		input_array[12][11][2]=41;
		input_array[13][11][2]=72;
		input_array[14][11][2]=55;
		input_array[15][11][2]=50;
		input_array[16][11][2]=64;
		input_array[17][11][2]=56;
		input_array[18][11][2]=69;
		input_array[19][11][2]=62;
		input_array[20][11][2]=43;
		input_array[21][11][2]=45;
		input_array[22][11][2]=61;
		input_array[23][11][2]=65;
		input_array[24][11][2]=68;
		input_array[25][11][2]=76;
		input_array[26][11][2]=79;
		input_array[27][11][2]=77;
		input_array[28][11][2]=48;
		input_array[29][11][2]=45;
		input_array[30][11][2]=48;
		input_array[31][11][2]=56;
		input_array[0][12][2]=48;
		input_array[1][12][2]=59;
		input_array[2][12][2]=64;
		input_array[3][12][2]=82;
		input_array[4][12][2]=61;
		input_array[5][12][2]=42;
		input_array[6][12][2]=33;
		input_array[7][12][2]=35;
		input_array[8][12][2]=47;
		input_array[9][12][2]=64;
		input_array[10][12][2]=50;
		input_array[11][12][2]=27;
		input_array[12][12][2]=35;
		input_array[13][12][2]=59;
		input_array[14][12][2]=57;
		input_array[15][12][2]=50;
		input_array[16][12][2]=47;
		input_array[17][12][2]=47;
		input_array[18][12][2]=50;
		input_array[19][12][2]=53;
		input_array[20][12][2]=58;
		input_array[21][12][2]=60;
		input_array[22][12][2]=58;
		input_array[23][12][2]=60;
		input_array[24][12][2]=56;
		input_array[25][12][2]=61;
		input_array[26][12][2]=57;
		input_array[27][12][2]=50;
		input_array[28][12][2]=45;
		input_array[29][12][2]=56;
		input_array[30][12][2]=56;
		input_array[31][12][2]=62;
		input_array[0][13][2]=70;
		input_array[1][13][2]=67;
		input_array[2][13][2]=84;
		input_array[3][13][2]=87;
		input_array[4][13][2]=78;
		input_array[5][13][2]=80;
		input_array[6][13][2]=17;
		input_array[7][13][2]=20;
		input_array[8][13][2]=36;
		input_array[9][13][2]=39;
		input_array[10][13][2]=47;
		input_array[11][13][2]=39;
		input_array[12][13][2]=30;
		input_array[13][13][2]=35;
		input_array[14][13][2]=49;
		input_array[15][13][2]=55;
		input_array[16][13][2]=64;
		input_array[17][13][2]=82;
		input_array[18][13][2]=97;
		input_array[19][13][2]=102;
		input_array[20][13][2]=93;
		input_array[21][13][2]=62;
		input_array[22][13][2]=66;
		input_array[23][13][2]=60;
		input_array[24][13][2]=50;
		input_array[25][13][2]=53;
		input_array[26][13][2]=55;
		input_array[27][13][2]=48;
		input_array[28][13][2]=52;
		input_array[29][13][2]=61;
		input_array[30][13][2]=56;
		input_array[31][13][2]=54;
		input_array[0][14][2]=68;
		input_array[1][14][2]=72;
		input_array[2][14][2]=86;
		input_array[3][14][2]=76;
		input_array[4][14][2]=77;
		input_array[5][14][2]=81;
		input_array[6][14][2]=19;
		input_array[7][14][2]=25;
		input_array[8][14][2]=36;
		input_array[9][14][2]=34;
		input_array[10][14][2]=72;
		input_array[11][14][2]=93;
		input_array[12][14][2]=81;
		input_array[13][14][2]=86;
		input_array[14][14][2]=97;
		input_array[15][14][2]=98;
		input_array[16][14][2]=71;
		input_array[17][14][2]=136;
		input_array[18][14][2]=162;
		input_array[19][14][2]=154;
		input_array[20][14][2]=133;
		input_array[21][14][2]=76;
		input_array[22][14][2]=65;
		input_array[23][14][2]=59;
		input_array[24][14][2]=65;
		input_array[25][14][2]=64;
		input_array[26][14][2]=61;
		input_array[27][14][2]=67;
		input_array[28][14][2]=54;
		input_array[29][14][2]=62;
		input_array[30][14][2]=48;
		input_array[31][14][2]=44;
		input_array[0][15][2]=40;
		input_array[1][15][2]=51;
		input_array[2][15][2]=61;
		input_array[3][15][2]=67;
		input_array[4][15][2]=62;
		input_array[5][15][2]=67;
		input_array[6][15][2]=32;
		input_array[7][15][2]=28;
		input_array[8][15][2]=53;
		input_array[9][15][2]=44;
		input_array[10][15][2]=99;
		input_array[11][15][2]=105;
		input_array[12][15][2]=102;
		input_array[13][15][2]=107;
		input_array[14][15][2]=112;
		input_array[15][15][2]=113;
		input_array[16][15][2]=85;
		input_array[17][15][2]=124;
		input_array[18][15][2]=153;
		input_array[19][15][2]=168;
		input_array[20][15][2]=145;
		input_array[21][15][2]=104;
		input_array[22][15][2]=90;
		input_array[23][15][2]=74;
		input_array[24][15][2]=78;
		input_array[25][15][2]=82;
		input_array[26][15][2]=77;
		input_array[27][15][2]=80;
		input_array[28][15][2]=61;
		input_array[29][15][2]=73;
		input_array[30][15][2]=55;
		input_array[31][15][2]=66;
		input_array[0][16][2]=33;
		input_array[1][16][2]=41;
		input_array[2][16][2]=48;
		input_array[3][16][2]=66;
		input_array[4][16][2]=58;
		input_array[5][16][2]=57;
		input_array[6][16][2]=61;
		input_array[7][16][2]=22;
		input_array[8][16][2]=54;
		input_array[9][16][2]=65;
		input_array[10][16][2]=116;
		input_array[11][16][2]=114;
		input_array[12][16][2]=114;
		input_array[13][16][2]=118;
		input_array[14][16][2]=126;
		input_array[15][16][2]=127;
		input_array[16][16][2]=109;
		input_array[17][16][2]=110;
		input_array[18][16][2]=131;
		input_array[19][16][2]=145;
		input_array[20][16][2]=146;
		input_array[21][16][2]=112;
		input_array[22][16][2]=103;
		input_array[23][16][2]=72;
		input_array[24][16][2]=73;
		input_array[25][16][2]=87;
		input_array[26][16][2]=88;
		input_array[27][16][2]=82;
		input_array[28][16][2]=71;
		input_array[29][16][2]=74;
		input_array[30][16][2]=61;
		input_array[31][16][2]=66;
		input_array[0][17][2]=38;
		input_array[1][17][2]=35;
		input_array[2][17][2]=47;
		input_array[3][17][2]=59;
		input_array[4][17][2]=60;
		input_array[5][17][2]=58;
		input_array[6][17][2]=52;
		input_array[7][17][2]=6;
		input_array[8][17][2]=40;
		input_array[9][17][2]=89;
		input_array[10][17][2]=117;
		input_array[11][17][2]=127;
		input_array[12][17][2]=136;
		input_array[13][17][2]=131;
		input_array[14][17][2]=125;
		input_array[15][17][2]=128;
		input_array[16][17][2]=122;
		input_array[17][17][2]=113;
		input_array[18][17][2]=113;
		input_array[19][17][2]=85;
		input_array[20][17][2]=115;
		input_array[21][17][2]=98;
		input_array[22][17][2]=77;
		input_array[23][17][2]=65;
		input_array[24][17][2]=78;
		input_array[25][17][2]=85;
		input_array[26][17][2]=93;
		input_array[27][17][2]=91;
		input_array[28][17][2]=74;
		input_array[29][17][2]=74;
		input_array[30][17][2]=77;
		input_array[31][17][2]=65;
		input_array[0][18][2]=62;
		input_array[1][18][2]=64;
		input_array[2][18][2]=70;
		input_array[3][18][2]=71;
		input_array[4][18][2]=65;
		input_array[5][18][2]=64;
		input_array[6][18][2]=54;
		input_array[7][18][2]=29;
		input_array[8][18][2]=49;
		input_array[9][18][2]=105;
		input_array[10][18][2]=120;
		input_array[11][18][2]=135;
		input_array[12][18][2]=145;
		input_array[13][18][2]=142;
		input_array[14][18][2]=127;
		input_array[15][18][2]=137;
		input_array[16][18][2]=133;
		input_array[17][18][2]=110;
		input_array[18][18][2]=100;
		input_array[19][18][2]=62;
		input_array[20][18][2]=77;
		input_array[21][18][2]=65;
		input_array[22][18][2]=53;
		input_array[23][18][2]=78;
		input_array[24][18][2]=83;
		input_array[25][18][2]=78;
		input_array[26][18][2]=88;
		input_array[27][18][2]=87;
		input_array[28][18][2]=79;
		input_array[29][18][2]=76;
		input_array[30][18][2]=81;
		input_array[31][18][2]=61;
		input_array[0][19][2]=64;
		input_array[1][19][2]=74;
		input_array[2][19][2]=76;
		input_array[3][19][2]=78;
		input_array[4][19][2]=64;
		input_array[5][19][2]=61;
		input_array[6][19][2]=68;
		input_array[7][19][2]=74;
		input_array[8][19][2]=73;
		input_array[9][19][2]=111;
		input_array[10][19][2]=126;
		input_array[11][19][2]=133;
		input_array[12][19][2]=137;
		input_array[13][19][2]=141;
		input_array[14][19][2]=132;
		input_array[15][19][2]=138;
		input_array[16][19][2]=137;
		input_array[17][19][2]=112;
		input_array[18][19][2]=61;
		input_array[19][19][2]=56;
		input_array[20][19][2]=66;
		input_array[21][19][2]=60;
		input_array[22][19][2]=58;
		input_array[23][19][2]=85;
		input_array[24][19][2]=86;
		input_array[25][19][2]=80;
		input_array[26][19][2]=79;
		input_array[27][19][2]=71;
		input_array[28][19][2]=77;
		input_array[29][19][2]=72;
		input_array[30][19][2]=68;
		input_array[31][19][2]=54;
		input_array[0][20][2]=60;
		input_array[1][20][2]=64;
		input_array[2][20][2]=74;
		input_array[3][20][2]=63;
		input_array[4][20][2]=58;
		input_array[5][20][2]=71;
		input_array[6][20][2]=77;
		input_array[7][20][2]=62;
		input_array[8][20][2]=61;
		input_array[9][20][2]=102;
		input_array[10][20][2]=128;
		input_array[11][20][2]=129;
		input_array[12][20][2]=134;
		input_array[13][20][2]=140;
		input_array[14][20][2]=125;
		input_array[15][20][2]=132;
		input_array[16][20][2]=125;
		input_array[17][20][2]=116;
		input_array[18][20][2]=36;
		input_array[19][20][2]=44;
		input_array[20][20][2]=51;
		input_array[21][20][2]=57;
		input_array[22][20][2]=60;
		input_array[23][20][2]=82;
		input_array[24][20][2]=76;
		input_array[25][20][2]=82;
		input_array[26][20][2]=73;
		input_array[27][20][2]=54;
		input_array[28][20][2]=57;
		input_array[29][20][2]=58;
		input_array[30][20][2]=55;
		input_array[31][20][2]=58;
		input_array[0][21][2]=44;
		input_array[1][21][2]=63;
		input_array[2][21][2]=64;
		input_array[3][21][2]=55;
		input_array[4][21][2]=73;
		input_array[5][21][2]=63;
		input_array[6][21][2]=61;
		input_array[7][21][2]=55;
		input_array[8][21][2]=55;
		input_array[9][21][2]=69;
		input_array[10][21][2]=100;
		input_array[11][21][2]=102;
		input_array[12][21][2]=128;
		input_array[13][21][2]=141;
		input_array[14][21][2]=122;
		input_array[15][21][2]=126;
		input_array[16][21][2]=116;
		input_array[17][21][2]=118;
		input_array[18][21][2]=21;
		input_array[19][21][2]=5;
		input_array[20][21][2]=30;
		input_array[21][21][2]=45;
		input_array[22][21][2]=59;
		input_array[23][21][2]=77;
		input_array[24][21][2]=61;
		input_array[25][21][2]=65;
		input_array[26][21][2]=57;
		input_array[27][21][2]=46;
		input_array[28][21][2]=48;
		input_array[29][21][2]=52;
		input_array[30][21][2]=48;
		input_array[31][21][2]=41;
		input_array[0][22][2]=18;
		input_array[1][22][2]=47;
		input_array[2][22][2]=38;
		input_array[3][22][2]=62;
		input_array[4][22][2]=66;
		input_array[5][22][2]=53;
		input_array[6][22][2]=52;
		input_array[7][22][2]=55;
		input_array[8][22][2]=49;
		input_array[9][22][2]=35;
		input_array[10][22][2]=72;
		input_array[11][22][2]=47;
		input_array[12][22][2]=64;
		input_array[13][22][2]=80;
		input_array[14][22][2]=44;
		input_array[15][22][2]=43;
		input_array[16][22][2]=100;
		input_array[17][22][2]=114;
		input_array[18][22][2]=34;
		input_array[19][22][2]=16;
		input_array[20][22][2]=14;
		input_array[21][22][2]=28;
		input_array[22][22][2]=48;
		input_array[23][22][2]=69;
		input_array[24][22][2]=50;
		input_array[25][22][2]=41;
		input_array[26][22][2]=48;
		input_array[27][22][2]=44;
		input_array[28][22][2]=50;
		input_array[29][22][2]=50;
		input_array[30][22][2]=33;
		input_array[31][22][2]=42;
		input_array[0][23][2]=17;
		input_array[1][23][2]=32;
		input_array[2][23][2]=40;
		input_array[3][23][2]=52;
		input_array[4][23][2]=56;
		input_array[5][23][2]=56;
		input_array[6][23][2]=46;
		input_array[7][23][2]=46;
		input_array[8][23][2]=37;
		input_array[9][23][2]=38;
		input_array[10][23][2]=62;
		input_array[11][23][2]=16;
		input_array[12][23][2]=26;
		input_array[13][23][2]=21;
		input_array[14][23][2]=19;
		input_array[15][23][2]=22;
		input_array[16][23][2]=69;
		input_array[17][23][2]=89;
		input_array[18][23][2]=39;
		input_array[19][23][2]=36;
		input_array[20][23][2]=12;
		input_array[21][23][2]=29;
		input_array[22][23][2]=27;
		input_array[23][23][2]=67;
		input_array[24][23][2]=51;
		input_array[25][23][2]=40;
		input_array[26][23][2]=35;
		input_array[27][23][2]=36;
		input_array[28][23][2]=35;
		input_array[29][23][2]=47;
		input_array[30][23][2]=32;
		input_array[31][23][2]=40;
		input_array[0][24][2]=37;
		input_array[1][24][2]=48;
		input_array[2][24][2]=52;
		input_array[3][24][2]=39;
		input_array[4][24][2]=49;
		input_array[5][24][2]=46;
		input_array[6][24][2]=43;
		input_array[7][24][2]=45;
		input_array[8][24][2]=43;
		input_array[9][24][2]=38;
		input_array[10][24][2]=49;
		input_array[11][24][2]=18;
		input_array[12][24][2]=42;
		input_array[13][24][2]=62;
		input_array[14][24][2]=58;
		input_array[15][24][2]=42;
		input_array[16][24][2]=48;
		input_array[17][24][2]=74;
		input_array[18][24][2]=35;
		input_array[19][24][2]=41;
		input_array[20][24][2]=29;
		input_array[21][24][2]=43;
		input_array[22][24][2]=29;
		input_array[23][24][2]=35;
		input_array[24][24][2]=65;
		input_array[25][24][2]=52;
		input_array[26][24][2]=44;
		input_array[27][24][2]=44;
		input_array[28][24][2]=31;
		input_array[29][24][2]=61;
		input_array[30][24][2]=53;
		input_array[31][24][2]=47;
		input_array[0][25][2]=27;
		input_array[1][25][2]=32;
		input_array[2][25][2]=54;
		input_array[3][25][2]=49;
		input_array[4][25][2]=43;
		input_array[5][25][2]=57;
		input_array[6][25][2]=54;
		input_array[7][25][2]=53;
		input_array[8][25][2]=51;
		input_array[9][25][2]=45;
		input_array[10][25][2]=46;
		input_array[11][25][2]=26;
		input_array[12][25][2]=54;
		input_array[13][25][2]=58;
		input_array[14][25][2]=54;
		input_array[15][25][2]=52;
		input_array[16][25][2]=57;
		input_array[17][25][2]=64;
		input_array[18][25][2]=66;
		input_array[19][25][2]=54;
		input_array[20][25][2]=32;
		input_array[21][25][2]=25;
		input_array[22][25][2]=62;
		input_array[23][25][2]=25;
		input_array[24][25][2]=62;
		input_array[25][25][2]=56;
		input_array[26][25][2]=34;
		input_array[27][25][2]=36;
		input_array[28][25][2]=41;
		input_array[29][25][2]=67;
		input_array[30][25][2]=51;
		input_array[31][25][2]=60;
		input_array[0][26][2]=37;
		input_array[1][26][2]=31;
		input_array[2][26][2]=49;
		input_array[3][26][2]=52;
		input_array[4][26][2]=49;
		input_array[5][26][2]=60;
		input_array[6][26][2]=59;
		input_array[7][26][2]=59;
		input_array[8][26][2]=57;
		input_array[9][26][2]=51;
		input_array[10][26][2]=46;
		input_array[11][26][2]=29;
		input_array[12][26][2]=60;
		input_array[13][26][2]=47;
		input_array[14][26][2]=56;
		input_array[15][26][2]=36;
		input_array[16][26][2]=49;
		input_array[17][26][2]=59;
		input_array[18][26][2]=73;
		input_array[19][26][2]=57;
		input_array[20][26][2]=47;
		input_array[21][26][2]=30;
		input_array[22][26][2]=67;
		input_array[23][26][2]=44;
		input_array[24][26][2]=48;
		input_array[25][26][2]=48;
		input_array[26][26][2]=34;
		input_array[27][26][2]=52;
		input_array[28][26][2]=61;
		input_array[29][26][2]=51;
		input_array[30][26][2]=31;
		input_array[31][26][2]=43;
		input_array[0][27][2]=43;
		input_array[1][27][2]=43;
		input_array[2][27][2]=42;
		input_array[3][27][2]=45;
		input_array[4][27][2]=51;
		input_array[5][27][2]=56;
		input_array[6][27][2]=59;
		input_array[7][27][2]=60;
		input_array[8][27][2]=75;
		input_array[9][27][2]=60;
		input_array[10][27][2]=45;
		input_array[11][27][2]=27;
		input_array[12][27][2]=52;
		input_array[13][27][2]=53;
		input_array[14][27][2]=56;
		input_array[15][27][2]=35;
		input_array[16][27][2]=29;
		input_array[17][27][2]=56;
		input_array[18][27][2]=51;
		input_array[19][27][2]=50;
		input_array[20][27][2]=50;
		input_array[21][27][2]=52;
		input_array[22][27][2]=37;
		input_array[23][27][2]=51;
		input_array[24][27][2]=56;
		input_array[25][27][2]=49;
		input_array[26][27][2]=60;
		input_array[27][27][2]=63;
		input_array[28][27][2]=58;
		input_array[29][27][2]=46;
		input_array[30][27][2]=47;
		input_array[31][27][2]=47;
		input_array[0][28][2]=45;
		input_array[1][28][2]=55;
		input_array[2][28][2]=52;
		input_array[3][28][2]=49;
		input_array[4][28][2]=52;
		input_array[5][28][2]=51;
		input_array[6][28][2]=50;
		input_array[7][28][2]=52;
		input_array[8][28][2]=63;
		input_array[9][28][2]=46;
		input_array[10][28][2]=42;
		input_array[11][28][2]=31;
		input_array[12][28][2]=48;
		input_array[13][28][2]=44;
		input_array[14][28][2]=37;
		input_array[15][28][2]=44;
		input_array[16][28][2]=51;
		input_array[17][28][2]=63;
		input_array[18][28][2]=47;
		input_array[19][28][2]=46;
		input_array[20][28][2]=52;
		input_array[21][28][2]=56;
		input_array[22][28][2]=46;
		input_array[23][28][2]=54;
		input_array[24][28][2]=77;
		input_array[25][28][2]=59;
		input_array[26][28][2]=57;
		input_array[27][28][2]=49;
		input_array[28][28][2]=46;
		input_array[29][28][2]=56;
		input_array[30][28][2]=57;
		input_array[31][28][2]=56;
		input_array[0][29][2]=52;
		input_array[1][29][2]=56;
		input_array[2][29][2]=52;
		input_array[3][29][2]=57;
		input_array[4][29][2]=45;
		input_array[5][29][2]=48;
		input_array[6][29][2]=55;
		input_array[7][29][2]=65;
		input_array[8][29][2]=72;
		input_array[9][29][2]=63;
		input_array[10][29][2]=47;
		input_array[11][29][2]=61;
		input_array[12][29][2]=58;
		input_array[13][29][2]=66;
		input_array[14][29][2]=72;
		input_array[15][29][2]=72;
		input_array[16][29][2]=65;
		input_array[17][29][2]=61;
		input_array[18][29][2]=58;
		input_array[19][29][2]=64;
		input_array[20][29][2]=64;
		input_array[21][29][2]=65;
		input_array[22][29][2]=68;
		input_array[23][29][2]=72;
		input_array[24][29][2]=82;
		input_array[25][29][2]=67;
		input_array[26][29][2]=60;
		input_array[27][29][2]=61;
		input_array[28][29][2]=67;
		input_array[29][29][2]=70;
		input_array[30][29][2]=61;
		input_array[31][29][2]=52;
		input_array[0][30][2]=51;
		input_array[1][30][2]=52;
		input_array[2][30][2]=56;
		input_array[3][30][2]=58;
		input_array[4][30][2]=47;
		input_array[5][30][2]=46;
		input_array[6][30][2]=60;
		input_array[7][30][2]=61;
		input_array[8][30][2]=61;
		input_array[9][30][2]=63;
		input_array[10][30][2]=59;
		input_array[11][30][2]=61;
		input_array[12][30][2]=68;
		input_array[13][30][2]=65;
		input_array[14][30][2]=82;
		input_array[15][30][2]=76;
		input_array[16][30][2]=62;
		input_array[17][30][2]=58;
		input_array[18][30][2]=62;
		input_array[19][30][2]=71;
		input_array[20][30][2]=61;
		input_array[21][30][2]=75;
		input_array[22][30][2]=71;
		input_array[23][30][2]=66;
		input_array[24][30][2]=77;
		input_array[25][30][2]=70;
		input_array[26][30][2]=68;
		input_array[27][30][2]=68;
		input_array[28][30][2]=66;
		input_array[29][30][2]=53;
		input_array[30][30][2]=49;
		input_array[31][30][2]=55;
		input_array[0][31][2]=56;
		input_array[1][31][2]=53;
		input_array[2][31][2]=53;
		input_array[3][31][2]=61;
		input_array[4][31][2]=61;
		input_array[5][31][2]=59;
		input_array[6][31][2]=61;
		input_array[7][31][2]=44;
		input_array[8][31][2]=40;
		input_array[9][31][2]=49;
		input_array[10][31][2]=53;
		input_array[11][31][2]=56;
		input_array[12][31][2]=58;
		input_array[13][31][2]=57;
		input_array[14][31][2]=62;
		input_array[15][31][2]=74;
		input_array[16][31][2]=62;
		input_array[17][31][2]=58;
		input_array[18][31][2]=55;
		input_array[19][31][2]=67;
		input_array[20][31][2]=54;
		input_array[21][31][2]=66;
		input_array[22][31][2]=53;
		input_array[23][31][2]=39;
		input_array[24][31][2]=59;
		input_array[25][31][2]=42;
		input_array[26][31][2]=44;
		input_array[27][31][2]=48;
		input_array[28][31][2]=38;
		input_array[29][31][2]=28;
		input_array[30][31][2]=37;
		input_array[31][31][2]=46;

        #20;
        reset=0;
        enable=1;
    end
   
    
    always #10 clock=~clock;
   
endmodule
